��   v��A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ����UI_CON�FIG_T  �x L$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�73�ODE�
4�CFOCA �5VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j �Ơ!BG�#�!hIN=SR$IO}7�PM�X_PKT�?$IHELP�� ME�#BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�<S�TYf2$Iv!_8Gv!k FKE�F�HTML�_N;AM�#DIMC4:1>]ABRIGH83s oDJ7CH92%!FEL0T_DEVICg1�&USTO_@ � t @A�R$@PIDD�BC��D*PAG� ?xhA�B�ISCREu�EF���GN�@�$FLAG�@�4&�1  h �	$PWD_ACGCES� MA�8��hS:1�%)$L�ABE� $T�z jHP�3�R�	>4SUSRVI 1  < `�R*��R��QPRI��m� t1�PTRIP��"m�$$CLA~SP ���a���R��R `\ SI��	g  �1N�$'2 ����R	 /,��?���aa1`jbed`a����� /� �`�o���
 ��(/SO�FTP�@/GEN��1?CURREN�T=>�A,952�,1 ���4/UUІ`��b�� 1 set �var ;g.`[?1] = '�o�`�  �o�o,378�,3�o�d�~2�/Ax)�_81,'10 w�bۏ~!3����}1����(s47�I�[��}2~����(s5��Axa _�q���������˟Z� ���%�7�I�؟m� �������ǯV���� �!�3�E�W��{��������ÿտ�� ?TPTX����l��� s ��鶄�$/sof�tpart/ge�nlink?he�lp=/md/t�pmenu.dg@޿xϊϜϮ�g�&C�U�pwdd����� 1�f�U�g�yߋߝ߯� >�������	��-�� ��c�u�������+�a�f�b�� ($R������6�!�Z���ada��c������� SW?IP[61]��dcH�g���aJ��aJ�  ��J�	H�������d���}�8�b���`  ���H �Gp�N�L#J�Ffbc �:c�B 1)hR� \��_}�� REG V�ED?���wh�olemod.h�tm�	singl��doub�tripbrows3b� i{�W������"/����dev.s�lo/� 1r,	t�/A�// K/�/�/?�/5?G?Y?8k?}?�?� ��? �?�?�?OO+O=OOOaOjE @�?�O�OpO �O�O�O�F�	�?�?_ /_A_S_e_w_�_�_�_ �_�_�_�_oo+o=o Ooao/'yoso�o�o�o �o�o�o1CU gy������ �? �2�D�V�h�z��� �����O���Ǐُ .�@��O	_������� ��П˟ݟ���%� 7�`�[�m�������� �oկϯ���!�3�E� W�i�{�������ÿտ �����/�A��|� �Ϡϲ���������� ��B�T�#�5ߊߜ� S�e�K��������,� '�9�K�t�o���� ����������߯1� +�Y�k�}��������� ������1CU gy��k����  2DVhzu� ��������� �@/;/M/_/�/�/�/ �/�/�/�/�/??%? 7?`?[?m?;��?�?�? �?�?�?�?O!O3OEO WOiO{O�O�O�O�O�O �O�O�4_F_X_j_|_ �_�_�_�_�_��_o��_�_BoTobj�$U�I_TOPMEN�U 1-`�a�R 
d��aQ)*def�ault_ ]�*level0 =*[	 �o�0��o�o�o	rtpi�o[23]�8tpst[1=xY��o�o�=h58�e01_l.pn�g��6menu15�y�p�q13�z�r��z�t4�{��q�� ?�f�x���������R T������1�C�҄�prim=�qp�age,1422,1J���������˟ ֏���%�7�I�ؖ�^�class,5R���������ϯڔf�13֯��0�hB�T�ۓ^�53p�@������ƿؿۓ^�8��%�7�I�[�ڟ�ϑϣϵ�����Y �`�a�o��mΙq�;�Y�CvtyN}6HqOmf[0PN�	�Пc[164=w��5�9=x�q)�o���x2 ��}Q����w�{�� O������� ��$� o�H�Z�l�~�����1� �������� ��e�22gy���> p���	-�� ��n����e�w�1���//*/</���^�ainedi�	�s/�/�/�/�/���config=s�ingle&^�wintpj��/??�*?<?����r?!ٙ�gl[57�ٕ�?$wޔ08�ݔ07�9�?h�6���62,O[6�:��?OqO�x��z�4s�x�O���x�  �B�Q�*_<_N_`_r_ �_���_�_�_�_�_o �_&o8oJo\ono�o�oz�!;�$doub�%�oc�13~�&du�al�i38��,4�o�o�o9�o�n�o �ax��#o��������%3.=_!g�Q�b8"�z��� ��U�\ԏ���
����+:6��i48,2�Q��b]������  ]?ҟ�/�UE��O����s��:�_���G�u �����n�l��O�J�h�M�;�6G�u7� �����ÿտ翦 ��/�A�S�e����π�ϭϿ��������"�1�/�A�S�e�w� �ϛ߭߿������߄� �+�=�O�a�s��� �������������6
�?�Q�c�u����$��74������������C���6�	TPTX[209�<aAY2+H,���BY1�8t?Ht���a
t0�2��aA��=�DtvB��O�L_��0��Li�S=�treeview�#�X�3��`�381,26�o//A/S/�w/ �/�/�/�/�/`/�/?�?+?=?O?�o���5��o%���?�?�?�ADr?>1`��?"2�� FOXOc?�?�_�.E-� �O�O�OxO��@�O0OC_U_g_��6�OF�'_ n_�_�_�_8�_���_ �S�_Qocouo$vo�o 핪o#�oS�o�o 1CUz�os� �����
��y� 3�Z�l�~��������/ ؏���� �2���V� h�z�������?�� ��
��.�@�ϟd�v� ��������M����� �*�<�˯N�r����� ����̿[����&� 8�J�ٿnπϒϤ϶� ��wo�o�ϭo"߉'� E�W�i�{ߎߟ߱��� 1�������/�A�S� e�w�9����������� ��e�>�P�b�t��� ��'��������� ��:L^p��� 5��� $� HZl~��1� ���/ /2/�V/ h/z/�/�/�/?/�/�/ �/
??.?����d?� �?�ߍ�?�?�?�?�? OO)O�?5O_OqO�O �O�O�O�O�O��_&_ 8_J_\_n_�_�/�_�_ �_�_�_�_�_"o4oFo Xojo|oo�o�o�o�o �o�o�o0BTf x������ ��,�>�P�b�t��� ��'���Ώ����� ��:�L�^�p�����C? U?ʟy?�UO�O�#� 5�G�Y�k�~������� ůׯ�����1�C� _z�������¿Կ� �
��.�@�R�d�� �ϚϬϾ�����q�� �*�<�N�`���rߖ� �ߺ���������&� 8�J�\�n��ߒ��� ������{���"�4�F� X�j�|�������������������*de�fault؞*level8a�໯Y�w�! tpst[1]�	��y�tpioG[23���u��d�,>men�u7_l.png�A^13cp5�x]�[4�u6 cp���	//-/?/ ��c/u/�/�/�/�/L/ �/�/??)?;?M?�"�prim=^p�age,74,1�R?�?�?�?�?�?�"�f6class,13�?OO0OBOTO�?�25ZO�O�O�O�O�O�#�<~O_$_6_H_Z_]?o218v?�_�_ �_�_�_�O�26�_o�-o?oQocoB�$U�I_USERVI�EW 1�����R 
���jo䒞o�o=m �o�o	-?�oc u���N��� ���o$�6�H���� ������ˏn���� %�7�I��m������ ��`�ԟ�X�!�3� E�W�i��������ï կx�����/�A�쟿*zoomT�?ZOOMIN�S� 񯺿̿޿�ϥ�&� 8�J�\�n�ϒϤ϶������<*maxr�esn�MAXRES���ω�R�d�v߈� ��=߾��������� *�<�N�`�r�߃�� ���������&�8� ��\�n�������G��� ��������3A ��|����g� �0B�fx ���Y���Q /,/>/P/b//�/�/ �/�/�/q/�/??(? :?�K?Y?k?�/�?�? �?�?�? O�?$O6OHO ZOlOO�O�O�O�O�O �?�O�O	_{OD_V_h_ z_�_/_�_�_�_�_�_ 
o�_.o@oRodovoa