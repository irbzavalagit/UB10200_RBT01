��   ��A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ����SEAL_M�AP_T  �0 �DI_��_�RDYT 8I�CFLTB	] QD�ISP>	wQFULLOPNB��	�CLS�	� �LT_STRB��QPRSSRRMB��Q� �BQH�I/Q( SEL8BNQVOL�
ko	ESTP	�o
8]�QCOM��QBUBL\	�o?RM1EMT~$�(2,."QMATbWBK$C)HIR)�HIC&TR_EMP_�%}(N�,�"})p��)�o
MOD
<� o	NSNG		1�	Wj'2'GH�(9C5QNOT_CaASc4�&0RA_��5�ART_OK���3QIN� OCB�4C'J\	�4C&�0��9�3c�7CQAUcTO�)5EC'NU�)�UEoEPRESE�'vD'UM+�CQ�� IN�0B�E�DETE�6�E})� \G|�D�ICHKP��U[Fn&5U�R_�ADV�VT�URGRQUE�vTmY�A}Y�A�HG_B�RSH��Ty8_BaYW�UQ�0E1BT�R�Z2�Z2�Z3�ZU3�Z4�Z4�Z5�Z55QG�NU�~gye�P_AC�3�gye�w)5�hye�X�fQA iwB�g�eK!�  u t{c2w�e�XPvKz�;viO_ONGU ��t�zd�u�z2d�u��zNd�u�zjd�u�z6�z6�wuQ|T/�)��x Q�)��xq�)��x��)� �x��)��у�u�P��톃u] ���uAB���EQ�u+��uSE!T(7G��ukC� `��uCL� ^��A�� p� P����uRLD�����G_W�0؛�u t�T�����v�A�) �Q;��uEND_JqO��]��uGOO_�{��ANE@�v��*��F��F��M��� ۥ�uw��u���vB�����;��uWAaIqn$W�#�DVTR82�z��vKTOuQ�v���}������uBLK8��ٵ�uUTH����ѶS���󩈙�7��h0A�h0)�INCH �y�q�V���A��X�� �ʪv}{-i�ű��vWi0���vsi�_I�#B�=�RAl�^�=��i��`v�c���c��MD�1� s�֩�ATM_AI�ש�w@�t����SSUR|S
��HAN��;t+��Sy���4�$$CLA�SS  ����r���!��!g�V�E+pONo��  1N�$�SLIO,  3 ~��! ��� �������������	� �D�V���z���w��� ��������
��q�B+Rs�(� �����  DV9z���� �_�
/-	/,
B,9/.