��   6��A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ����SEAL_S�CH_T  �� COMME�NT 'A�MOU= AT�OM_AIRNE�Q_ADD_DE�LAYN EQU�IPdGUNON�sFFdC_FA�CTOYC_BI{ASNPRE_� _S_TIMjD�=EjRAMPjR��i��xS_U�SEDN DUM�MY� HORMܲ �SUR�FLOW_TYP��%MOe jS�_wOFSMSEBwRSMGFSEM2G	2)n^ en�b	n�	��GUM�_DROP�4��$$CLASS  ������� �� �VER�SION��  1N�$�SL, ED1 3� �  d �1��=/��?�E/��  m(t'j/V*+/�/�/ �/s/�/�/�/:?�/^? �/b??'?�?K?�?o? �?�?�?6O�?ZO�?�? O#O�OGO�O�O}O�O �O2_D_�O_�Ok__ �_�_U_�_y_�_�_.o @o�_o�_goo�o�o �o�ouo�o�o�o< `�ocO)�M� q���8��\�� ��%���I�ڏm�� ����4�ǏE����� !���ğW���{�럟� 0�B�՟	���i���� ��S���w�篛�,�>� ����e�Q�+����� �s��Ͽ��:�Ϳ^� �b��'ϸ�K���o� �ϓϥ�6���Z����� �#ߴ�G��ߍ�}ߏ� ��2�D������k�� ����U��y����.� @������g������ ����u�������<�`��cO) Us�ed in MO?V_SEAM�� �s��):�^ �b'�K�o ���6/�Z/�� /#/�/G/�/�/}/�/ �/2?D?�/?�/k?? �?�?U?�?y?�?�?.O @O�?O�?gOO�O�O �O�OuO�O�O�O<__ `_�Oc_O_)_�_M_�_ q_�_�_�_8o�_\o�_ oo%o�oIo�omoo �o�o4�oE�o !��W�{�� 0�B��	��i���� ��S���w�珛�,�>� ����e�Q�+����� ��s��ϟ��:�͟^� �b��'���K�ܯo� ������6�ɯZ���� �#���G�ſ��}��� ��2�D�׿���k�� ����Uω�y��ϝ�.� @������g�߬߾� �߅�u����߫�<�� `���c�O�)��M��� q�����8���\��� ��%���I���m�� ����4��E�� !��W�{�� 0B�	�i� �S�w��,/>/ //�e/Q/+/�/�/ �/s/�/�/�/:?�/^? �/b??'?�?K?�?o? �?�?�?6O�?ZO�?�? O#O�OGO�O�O}O�O �O2_D_�O_�Ok__ �_�_U_�_y_�_�_.o @o�_o�_goo�o�o �o�ouo�o�o�o< `�ocO)�M� q���8��\�� ��%���I�ڏm�� ����4�ǏE����� !���ğW���{�럟� 0�B�՟	���i���� ��S���w�篛�,�>� ����e�Q�+����� �s��Ͽ��:�Ϳ^� �b��'ϸ�K���o� �ϓϥ�6���Z����� �#ߴ�G��ߍ�}ߏ� ��2�D������k�� ����U��y����.� @������g������ ����u�������< `��cO)�M� q���8�\� %�I�m ��4/�E//�/ !/�/�/W/�/{/�/�/ 0?B?�/	?�/i??�?��?S?�?w?�?�=�$�SLSCHED2 3 ���8A_ �0��?�ZOO~O�?�OmO)H3 5OGO�OkO_�O_�O'J4�O�O�_	_�_-_�_Q_'J5q_�_2o�_ Vo�_Zo�_Ca