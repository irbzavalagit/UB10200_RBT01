��   #�A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ����CELL_G�RP_T   �� $'FRA�ME $M�OUNT_LOC�CCF_METH�OD  $C�PY_SRC_I�DX_PLATF?RM_OFSCt�DIM_ $BA{SE{ FSETC���AUX_OR�DER   ��XYZ_MAgP �� ��LENGTH�T�TCH_GP_M�~ a AUTORA�IL_4�$$�CLASS  O�����D���DVERSIO�N  �1N�8LOO�R G��DD<Z$?���q���M,  1 <D? X< [�����Dk��i�����iO/�a/s/A/�/�/�/$ �/�/�/},�/0?�???m?7/�/ �?�?/�?�?	O�/!O�3OEO_I�$MNU�>A�2��  � <i�7���캷�?��ʺ7�;� "e� 2Ǻ���k�@�EZy��E�� đ���iy?�O��O_ �O_-_[_A_c_�_w_ �_�_�_�_�_o�_o Eo+o�O�O�O7oYo�o 1o�o�o�o�o/' Iw]���� ���+��3�a�G��Y���}���8�=�����ڀՁ����) ��O,���D��Oe?����Ď�q�=���U�Ï]��� q�����ӟ��۟	�� �?�%�7�Y���m��� ����ů�ٯ��;� !�C�q�W�y������� �����AX0ݿ�� U3�[�A�S�uϣω� ���Ͽ�������)� W�=�_ߍ�s߅��ߩ� ��������A�'�9� w�]�o�������� ����+��#�E�s�Y� {��������������� '/]CU�y ������	 G-?a�u�� �����/C/)/ K/y/_/q/�/�/�/�/ �/�/�/-??%?c?I?�  sGNUM  m�  �D v`��3TOOL}O�K��;�.�v0v1�13��0���.3�0������1��1'�ĈS3D?%� A�{?+OϿ3OaOGOYO {O�O�O�O�O�O�O_ �O_/_]_C_e_�_y_��_�_�_�;��?E*_ĈT<D�_�_ Jo�_Ro�ofoxo�o�o �o�o�o�o4, jPb����� �����8�f�L� n�������ҏ��ʏ� � �"�P�6�H���l� ~���Ο��֟���� :� �2�T���h����� �� ob�1a'O2j �o��ɯs�S?{� ������ÿ�׿��'� �/�]�C�U�wϥϋ� �����������	�+� Y�?�aߏ�uߗ��߫� ��������C�)�K� y�_�q��������� ����-��%�G�u�[� }��������������� )1_Eg�{ ������ I/Ac�w�� �����/E/+/ M/{/a/�/�/�?�4�3 �0�?