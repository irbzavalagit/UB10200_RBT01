��   4�A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ���	�SLGN_S�ETUP_T � H HPRO�C_WET_RU�N  UIF�_CYCLE_T�IF JLAST�MVGUN_ON�1 W	n VVOLU�MEV
� VSEA�L_AMO �YATOM_AI�RVPRESSU�R1�2VPAR�T_IDF JOB_ST�T�n^�:�n ����E��e�� � S ��S�CHEDUQ NU�M�TASK�FINIS�F�C �NINGFSLS�.WIZ� SL�CSTM_CTR���LOe�T�PP�BFRCA�LL��G�DS�B_AP_# FD�EFAULT_A�C�JNTWAR�N_EN,"USE�NONE4MAI�E� _F6 INT�F�MAJb*SEQ_IMPv*_!g%�RECOV�OKn|760�AD��MCSD�,REF�C��"S� Ef!4��*5�*6�*7�*8�*9�*10-;�08��083-;�+1�+1�;1;1;1,;2;8R� ��7��7h1��8�!�8�!�4SHO�RT�!H�0DU/BYTE�AH��PIh1PI�!& PL�_R_EL11� @ I��"A?TA_TYPk�B�INDEX�VA5R� R�=�$J2+4�G21�O�O��O�O+$ R�� f!_ARY �3 ;Q�1BT� PL, SPR_R0�^X�_W�2 ^XB^XB^X1mY1 mY1mY,1mX:2�Yi\ X2�Y�\v2�Y�\�2�Y@�\�2�Y�\�2mWIhR�hY2�hh2�h�"�h �"�h2�h2�h2�h ,2�g:3.x�lX3.x�l v3.x�l�3.x	|�3.x()|�3^VBhR�x� �yh1�y�!�y�!�y1 �y1�y1�y,1�x:2 m��|X2m�	�v2m�)� �2m�I��2m�i��2�wShQ%�� ,�h0 ,�� ,�� ,�0,�0 ,�0,�,0,�:1��)� X1��I�v1��i��1������1�����1%���,T �P�OSSIBQ OP�T }!LECT�EDz�� EQUI�0 �DM_FACT�O�IDQ FLO�WCM���_BIASV� ��� ��oPURG�0AT���n ǡ0Ih1PU_P�DTH|�!�>k#X_WAI�#ISP_SIG;��_!C�ån T� Y�2�Z�S�"R�����_�Cj"HI�*�L�O��VC3�����INù4��̳�3�� �α��������� �k"�9���29�XŮC�MOD�c�L�N_
 y�TMOU�_!��GRAVI�TEP C�+�_!Sࡨ4ą����_CNpu���â�_SQ� �  ġ
��L0Y!�)֢�A2(�F� ���3���3���3��C ��C���R���R���R ���Rb��Rb�j�cb� ��8cY�j�ġw�ġ�� ġ��ġ��ġ��ġ ��ġ������#���0�9�8c
 2P@PH$���SPEED1i_����2��NOΰ�a�P��R )�EPA �R������2��B���W���A��O�G�Ŏ_��VHOȄ: Q%飚�SAMPQ ����
 ���_O -AF^�S_D0S -A3��_N{��N�LOO�����BER��CON�Vc�)+�IO_C�OU��LDBGF�L�X�cRC_D�ELA��BRA�KEu�OVRL~"TBF_OFS	T`�S^��kO �MOPGGC�URR�Zz�AU�TO_�_T{F�DU����FZ �%̡AN � ��PcRP. �.OC6�|u�q OC_LA�mO�REe�THG �A��{ �T1V�A`w������SM� FP���H _����<O �DJDL��
 4����������������%����SEC�D���PR��BI J�cZ&2�Z&�2Z&B�Z%2c*2q*2*2R�x�2��%`�����!Hw1F�d�62�6 �26R�	5B6�R6 �R6�R6�R7�R7 ;c7-;8cF���4 55��4�9I5V��4e5 l��4�5���5�9�6�� �5;4����~CĥڣA ָ2��5?LPu�F�7���Ey��DRM�T�@�����BU�BT���� _OL�D_IS��)REQ� ��C��_ST=A��  IQW��9"TYPPRB;�CcOM��DU+ЉU ���@�XN�U�� �$� N�� �#��m�VYr�Vir�V yr�V�r�V�r�V�r�V�r�#R`�j�Efw��'�j��2��UBYTEj��h2�iiq�i�yq�4�SL�PL_P_��i� \ J��� g86���RAM�e�b 3s |Yswir�cQQi��� _�aLAz�R��3 ���_NA��%EX�JP+�FAUL��BOOKMARK��N��TCPF�LS"】w����x�v�?RTD�P�s�w����D���u�w���x���MQBIT�m*�f��w���K����AVG��TOe�������� C��_m���R���R���b��bIQJa�� ��2���B�������I2N�TR�R0T�@�2� ?�B�?���?�:�W2?� e2?�s2?��2?���Ϙ�J���Ϙj��Ϙ:�1���1��1��1ʜ2ڛII��Q��s���R �b�b�#b�1b �?b��1������� �������ʬ9��@�Y��
�y���BI����aιB�ι�aι I1ιW1ιe1ιs1ι�1θ��ηSI���`� �`m�B�mʽ`m�I0m� W0m�e0m�s0mʁ0m����%�b6�:u g� 	�pMQON  q<PLR�t����%����Q_E8�$�U��wU7�o�rv?�ATU�DP���`USR�C� � �� CUSX��AFLOW_CMN�{FL��D_TY����ID���н�ACC�����S �����IN�@�Кs�� %���2��Q-��7�ND�}�5��P�D�Й���հ����_ �_�_BoTo�B���"   �$$Cp�S  ����L�>�>� A�V�ERSIONI��  1No�$SL� EQI�l>�u� r���{�EQ
!��X�q��7GNS�Q3 j����,����>��*����	-9�SLWIZARD9f�����������>��@�R3~���  �s>�C>�)?��(@}�{d  ����2�^A jE�� C�^� ��� =��������/// �(H%�H)H/f'/ �/�/>/l/b/t/�/? !?�/�/<?"?{?�?s��>��,�?n(MOV_HOlp �?�8�3Q�?�?Р�7OEJ@ @>���CH!m@  �S�EH{���EO C ��?�O�O�I
w�B�3~�?�1>��34PNT�O;_2 �<P]0?B?�_b_�_�_p�?n�_q �/�,k�>���Я  '�P,i= ,oro�o�oYo�o�o�o �o&8�o\n �C����So� 
��.��R�d�v�9� ������Џ����� ۏ<�N�`�r������� ��̟ޟ���&�8�J�V�%V�z�e����� ¯���ѯ
���@� +�d�O���s������� �Ϳ��*��N�9� rτ�oϨϓ��Ϸ��� �����&�J�5�n��L��ߡ߳��TATUoS 3������ ���-�?� Q�c�u������� ������)�;�M�_� q�����������T�wL ��/ASew ������� +=R�as^� �����/�'/ 9/$/]/H/�/l/�/�/��/�/��USRCSoT 3�� X�&�ie"?4:H?��V�OLSET1  =�G�O���a:I2o?b93�?b94�?b95�?  