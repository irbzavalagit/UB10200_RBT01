��   ?3�A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ����MN_MCR�_TABLE �  � $MA�CRO_NAME� %$PRO�G@EPT_IN�DEX  $OPEN_IDa�ASSIGN_T�YPD  qk$MON_NO}�PREV_SUB�y a $USER�_WORK���_�L� MS�*RT�N  4&S�OP_T  �� $�EMG�O��RESE�T�MOT|�H�OLl�� 2��STAR PD�I8G9GAGBzGC�TPDS��REL�&U�s �� �EST�x��SFSP�C���C�C�NB��S)*$8�*$3%)4%)5%)6�%)7%)S�PNS�TRz�"D�  ��$$CLr   O����!������ VERSIO�N�(  �1N�:LDUOIMT 3��� �����$MAXDSRI� ��5
�$�.2 �%� � d%C�LR OF TR?ANSFER����%  L, U0a?���" ��q2�?�?�? �?�9���?!O�?EO�?�O{O*O�O�O`OrC�MOVE TO "�Ol5�@#_��KX���6tA�EREPAI[?l7P�IPN_�O�=	AT �POUNC_�KA�T�_�_�_%�f � MP EA�RLY�_o4PNC�LMZ?�_�_IPOS�IT� cEoo4na_�CL�oKo�<�EPURG�__[�a�o�o��]DISg SE COMPL� Ep3NDJOBI�? �����O��� (���#�p����C� U�ʏy�� ����6� �Z�	����?���Ɵ�u���DEFAU?LT ACCɟ�j#F_��˟�}��c�Ю���ҟ��! I�/O��g:!_I����\�-V��M�E?CHO OPsa����H�"�'�[FA�%
�STY1 ��:������Z sF��  �PATH���K� _��^[ѿ%WA?IT NEX��KI�S�^^5�{���w� �ϛ������:�L����5߂�1ߦ�U�g�T�urn Tabl�e Move T�o Pos�� TP�Ao`�߸���k��ENTER FIXT-ZON��=�NTRC�Q�Zx�:�EXK�C�T��i�Z^J��%=�I��BV�R�^0���� ����p�^KU��� ���� ��i�6��Z�l�aCLO;pV�AL�@1ml8SV�1T�q/T��2���
2����
3�5�
3&8J�
4���
4����
5���
5� //�
6�a/�
6R/d/v/�
7��/�
7�/�/�/�
8�)?�
8?,?>?�
9D�?�
9~?�?�?�
	0�?�	0�?�?OUO �OT�OxrO�O�O_��O�O�	b��OPN �_hOB[b\%�_ �_CZib\��_�_CZ �b\�Ko]oCZ1/b\ Q/�o�oCZ�/b\�/ %CZ�/b\?w�CZ ]?b\}?��CZ�?b\�??�Q�%EY&Oc\ EO�����=�_a�(_�"���F���j�|���V�ACUUM CAgN1 &���ACqP�џO��2 ���Pe�5�G���3d��9`ɯ������4ȯ��`-������5,��p��a�s���6���ep��ſ׿��7����pY�)�;���8X��-��ύϟ���9�����(!������0 �� ����V��������� ڟ��I���m��.�x� OFF}����� h�Z���x�����ﾩ 8�ܭz�J�\�"���@� �������� ��B $�dͦv�N� �l�
����,�� n>Pِ4����y����7//�� �/�/�/�/��/�/�/x?�/3_BLOWX  ��2NX0q_0?z/T5�n?OF�_�?�?T5w��?OF9o�?
OT5��6OOF�o\OnOT5?�OOF�O�O�E��OOFe$_6_�Eb_OF��_�_�Ek�_OF-��_�_�E�F*oOF��PoboU5 4/�o�`�o�o|/=O :s:?4�X�| ����9���o� ���B�T���ۏ���� ����5��Y�k��,� ��P�şt���������1����Rec P�ath Star�t5��dAERE�CSTAq��i	��b�Z�Pausse��}�PAUկڟ��%]�Re�sumί}�RES�9�����%]�Esnda�{�END������u�%Do Bwd Exij���h	DOBWDE'XITϠ��ٿ� `����?�ퟺ�i��� �ϟ���&���J�����
Sen�vent����S��EVN϶�j�=�%	}�Dgata�ߘ�DA��ڽ����%}�Sy�sVar��SY�SVY��(s��G�et��Z�GET����cz�quest Menu��~��REQMEN���첣��Prom�pt Box Y�NI�|�PROMP�T|����]�Y�q�M3sg����OK����=���%	Li�L?%LIST8�����%C�tatus�=]�TATPAG�E����%O;p.��try���OOPERe�����%Clear /User`�g3���USERCLRy����]�%For�cej������� �?�</;�`/_�ߖ/ E/�/�/{/�/?�/&? �/�/\??�?�?A?S? �?w?�?�?�?"O4OO XOOO�O=O�OaOsO �O�O�O_�O�OT__�x_'_9_%	Gri�p`�i���GRIPgPAR���jL/̇�fse�_��DR�O�_�_�z�a P�res����CHK�AoRo��b�Chec�k Noo���`N�OP�o�\C�o%~~`pare t�`�ick"KTO�PIC�[Y-%�eIqrocee���nULR2PRC踿�_��Z�Tur�n ON Vac�uum�}�VACOUUMO���[]�%	�FF�#�5�iF���Z\Y�%m�Blowoff����BLOWr���[�B��%S��Cu{rr�`Valv�~nUETVALV���4��MH To�olq�R�_TOO  c͟|�"/�f_'�֟ �_"�o����B�T�ɯ x��������5��Y� ����>���ſt��� �����ο�U�g�R� ��:�L���p��ϔϦ��BYPASS ROBOTq�����Pқ���������v}$�AUTO ӠY�@�8�^�pӖ�u��$MACRO_M�AX/����0���S)N�BL �����՗�b�b�A���>�PDIMSpp��f��Y�SUc��u�TPDSBEX�  -�q�U� �������