��  	�A��*SYST�EM*��V9.3�0126 2/�12/2021 A�  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ��4�AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�>#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@!LRM_RE�CO"  � A�LM�"ENB���&ON�!� MDG�/ 0 $DEBUG1A�"d
�$3AO� ."��!�_IF� � 
$ENABL@QC#� P dC#U5K�!MA�B �"��
� OG�f 0COURR_D1P $Q3GLIN@S1I4$C$�AUSOd�APPINFOEQ/ � �L A �?1�5�1 H ��79EQUI�P 3�0NA�M� ��2_OV�R�$VERS�I� �!PCOU�PLE,   �$�!PPV1CES�0�!H  "P�R0�2	 � �$SOFT�T_�IDBTOTAL�_EQ� Q1]@N�O`BU SPI_I�NDE]uEXBS�CREEN_�4nBSIG�0O|%KW@PK_FI0�	$THKY��GPANEhD ~� DUMMY1d��D�!U4 Q!R�G1R�
 � /$TIT1d �� � 7Td7T� 7TP7TU55V65V75V85V95W05W>W�A7URW�Q7UfW1pW1zW1ʄW1�W2�R!SBoN_CF�!�0$!J� ; 
2�1�_CMNT�$�FLAGS]�C�HE"$Nb_O�PT�2 � ELL�SETUP � `�0HO�0 P�RZ1%{cMACR=O�bREPR�hD0�D+t@��b{�eH-M MN�B
1��UTOB U��0 9DE7VIC4STI�0�A� P@13��`BQd�f"VAL�#ISP�_UNI�#p_D�Ov7IyFR_F �@K%D13�;A�c��C_WA?t�a�zO�FF_@N�DEL�xLF0q�A�qr�?q�p�C?��`�A�E�C#�s�ATiB�t���bEX
 ~�! � 7( AX_y� x@-q�2qH�^`�1QrXu!P�EE�h�/0TOT��RE�se�^��b<�i�_RDYR&���IA �GW. 8 K�;@d�K�&U�eA�CB�� ��D"; . ?'� )b�C"SCAN=�g�=t�PO%Q� D� AVAIL Iq�l�Ҁ��r������� �, \�����A�!RDINqG�Bi�ԕCOM@�Tq��A�CSԗPI�R�AE� ADY��"MO� �sE 	� [M�s��2�REV�Bo�G��1�XI� %�R � � OD}`j�_$NO`M�C!b�x�/�"�u�� �������@D�d p E R�D_i�{ � FS�SB�&W`KBD_�SE2uAG���2B "_��B�� V�tp:5`סQC  ��a�_EDu 0  �S C2��`S�p��4%$l �t$O�P�@QB�q�_OqKࢃ0, P_C� �y��dh�U �`LACEI�!�a��֑Err�M� �0$D���֑�@�pX��OR BIGALLOW�G (KD2�2�@�VAR5�d!��L8[@S � ,KJq��H`S�pZ@M_Ox]zŗ�CFd7 X�0GR@�=M�NFLI����;@U��&�$� SWIT=$=�No`Ȓ��u_�G� �0WARNMxp�d��%`LI�V`NST� А-rFLT�R�TRA`�_T|�`� $ACCq�S�� X�r$OR�I�.&��RT�`_sSFg�CHGV0I�p�T�PA�I��T�A���� � �#@a�N�HDR���2�B�J; �C��3�4��5�6�7�8��9�!e`��x@�2w @� TRQ���$%f��֠����_�U�СᬐCOc <� �϶���3��2��LLEC_�>-�MULTIV4�"�$��A
2FS��IL�DD�
1��Oz@T_>1b   4� ,�6�1�=@�)24��x�0D�c! |9 $��.p��6�I`�L* \�TO��E��EX{����הI�� 2 ���"�@1�1b.'�����G�Q� #�"Q�/% �a��X�%�?sQD�UA$S�2�;A���M�� # C�NPO�% L�0a$# �X��pA��$JOB`B�Ъ����IGO�& dӠ��X��-'x��G�� �_M���' tӠF�L<�BNG�AW�TBA� ֑�!��/1��à�0���R0+P`/p%���`��(
Ё|��BqF!]�
2J�]�_RN�U�C`,J�`�e(�,J?�D/5C��)�����@V���P�_�`O3��a)��a$���8����IT�s��NOM@�3�c 2X����5TU�@P]�V�� ��*+P���� b��P�)����RAM��<��0�2A�z�
$TF32��D3
0����SU�`�!}�)m1H��p1�:EC��������A��Q��Ql3Y�NT>P��PDBG�DE'�+D��P����qt���+���AX��³uTn�AsUFpۦ��?AU1, ���lPFV`PI+�+m0P�GM�HM�IB@�F�F�GSIMQST}O�q$KEESPAT��z�28B�3hB���C�-S��0��`JB����aD�K�hY� gU�����. �U�CHNS�_EMP��$G��0�W�_�0�c;�1g_FP)5�0TC�Vn�T1�`%��T��%aaV����W"��JR��~��SEGFRAq��b��RST��LI9N�KcPVF��R�1CC/����kbZ"���Pbzr�"5(0` +�/��EՍa�P� �adP��Ar�d���idQ�SIZh��	t�fT��c�0z1y�aR��F �![�cP`'�ic|1`cx�P<`L���0�P�vCRC����]Ѓ �u�1`�x�Q���R�MI�N�w�Q`!�x�q�uD�����C��� ���`K�ݠ��R�EVR�� �Fh�_	eF�PN@��"�dQ�&��;�<�5�jc /�1V�I�|�0A��g��1� 1) a� SFV$�p#�1b���#�0�42= 2�Ќ�?��RG���"a�F@`���QqDcq��PLEW�!-�r�p<�ď֌��Rɤ3����������� U��R� HA;NC��$LG5б�@��Ӱ]@٠F���Ae���3�PR���S@���0��@�@@;�RA��@�CAZ�P��N��5O��GFCT�ѩ���F��p�r�PPPb ADI�O�a��a��&�Ӥ5�5����S[�g!�N�BMPUd(pY3�Q�AESpj���W��N  ShXYOZWPR�����⇶	/!�В�4 � �pI84��!5��n`_C�DϱW#�hN0'���6K@$��YC����&�SFLG������v�"-T(�[A��;A'�~�7� 6$��SUPp�ARM ����'��P]@8A� ��A��KP�#��x���UO��O��F��F���N��N���%n�GRqV~�O�'�DKI��sDK+3:�SUL���Vҷ�DD3r�GA*��R?�RK�RWܩ�
��Rw�R���:.�OOR��U>`�  ���ԯQ� q�:1��1打UTOOL �K��K��K�*�K� 7�K≓�¸���㊰�U��V��*���X��U��Y��Z��NU
��V��W��$�����<�E����URS�CC�T 8 H����`�� ��P_I��sL�k�k�d�IDX�1��2��3c��C}UPMMENU�]9)TITU����G%E!Ca:BZ_�#��: ��0�$ ��AS��&NO_HEADE��b��m��، �P�r�sx��T.��r�83��; TA����IRTR�P�w�x�L��,�C�0�RJ��t4��AERRL����<�"&q� OR��b$�j�`�00U�N_O7��P$S�YS� T � k�� 1�V�3V`B�D�BPXWOA�V0=�`$SKo1�BM]T��TRLU1>����pN`�4[�IND�ppDJ�$LAY_���A����PL��a_RWA���E?SERVED����A%r�"�UMM3Y9�10ِ�DB��U1?^�AP�R�q�P�DPOsS_�@U1@ ��������L7)ALD/�q��pV0Bj/�V#PCU1C�/�ql_�PENE�0TN��D�/@� REC|��U1EH m0�O�`@$L�#A$7#�B{�;R`�aUb�_D��@ROSSUbT�j��� �Ι@RIG6\6PA�USZ3TdETUR�NZ2�sMR_�0T�UC0�q)0EWM|Db"�IGNAL)���B$LA\�5f�B$P,�C$P̬�ހD�0��PC�4���pDO^`,�&2�1�r*6GO_AWAY:2MOBa
¬B��DCSSҰST�CY_ F L�� �0�P��TB��]E2*XJ2fFN@O��|2躱@Bv�I50 G3 P����RB�b-��PIfGPO�HI_#BY���C�GTVr?C�HNDG�"HU���C�C�P�DSBLIOL�0TgF)�֖>DLS�QIR��O�UTEYFBt\m�FE41�֘SgD?C�bű�J��DOU��"�MCS�VbP(�R�R!r�HɠWİ�D.@M�SELE�L�T[`�Q�K� $w0��INK_NVsGb��b���FHA[Fq{p$
< Ayr"AA�A�wL ��MDL0b 3K��NR\��r��ce���j�c�e�cJ �c{r�de���mtw�P��}p�b��4!AA�SLAV�"M  ̰INPrP�FqPeyX?A����N�C� \��:   bL�wyX!�sSHOW�O 4���@�a�q�ra�r�v�u�v�r~��P` ,$\� r�����V���bS��:�ID������Wx�D�NT�V£�VEԴ�S�KI��遹S����2$D�QJ��;�_� Ǆ�SAFcڇ_SV>l�EXCLU����ONL� �Y�T1�ȠeHI_V��]�PPLY�R�y�HI`�0�_M�В��VRFY_d�.�M����OC+ Oճ��� 1D�����O�@3�LS��N�$e4���gC$`�_TPF$ED��Ab�CN��N���gEݓ8�@ճ�CHD0�0Qa_0e܀4PCPe���T��/ NB_V�AL���u�qQ 3Q� aTA�°N:  <DK`Cb R^rM�0j0��d����N?C'c"�S D $FP�_x�Fc�!I0p�_���H��~uA�PK_ T<��)�MARG��Ϣn�`S ~uSGO�U ���I�0�1 �18�j�< ��0An�|A~�ANNUN� @���gEI�d�0� ƹñ� ˺�YRE�F� I�!V @�> F����	$TOT�0�C$��$Ǔ��l5 EM�@NI�aCWOBU�)U�A���s�DAY�LOA�D�D�N��5"�EFF_AXIcR%X� �5�O��@�*�_� Q{Y٠O (��,r��E3����� 2X��(P�8�����D�A ��{Z 0�2чc p(2�C��K:SU�0W��E�yCA4p [��3 � �`�0IDLB5�W��-�+��V�G�V_-�й �DI�AG��{\� �1$d�`!�TAC �/q��'Q�����.r�R�"��,tV
 ��SW�1�Ђ�Ȁ2���Y0p��OH���J�PP
.rIR��.rBW��s��2 -q�~��w�/�0�x��Fn��[�������oRQDWg�MS` ���A2 O��,tLI�FE����!;rN@���#�ñ���CQW�³C9@�/@N�0Y����1FLA.�ñO�V90/� �0.rSU'PPO� �;r�1_��t�R�_X!2��)A��Z��W��9A��0&��"R!2XZ�q,t+Y2C9 TAB0B��NY���ñr _��-r�rICT��] `�PCACH����~ycv���2Nޕ�UFFI��@��Gq����6�CSF�DMSW�p^ 8۠KEYoIMAG3TM1�o��J��crJ=AO�CVIE$��_ �aBGL~�ð;��?� 	ǡu��`�٠�PST��! d�lǐl�pl��lEMAI�`V1[��5 5�FAUL]�a 4U3[�U�5@U���LTT6� bD�Pf�I������ ���=P�Mc�!���I,5�YRT� �Qc�< $N#�US�-Ў�IT9SBUF��;���DN��SUBz$�DC:�<QO"f�"SAV�%�"��@5r1.��'�ǶP�$N�UORD%�4�_z ��%`�"8OTTf�_5�[�Pm�MG�K4��FH7AX�#�x�Xz ���#_G�LqYN9_o�d <����ѕD�En�MY�*i�TϐF�>a��D5!�EDT_HP ��/e^r$�G�!"�&h�S`d����P�z�F5P f (�pSV^ �D���1��~qAФg� �����)3C_R/IK'�pB�mDVp�R�lE�ADSPdPBP�`�IIM�# �C�A<�Ad�U�G��4nCM�IP�PCX�T �DTH4 �S�B2��T2�CHS�3�CGBSC��C ��V�d�^VXP�#`T_DMcCONV�GMc`T4 $�Fz F�;pd�C�0�o1(�SC��gebCM�ER)�AFBCM�P)�@ETc mh�FU��DUn b��7�CD�Ix*P<0��EOӰB�i��j�XQ(�Q��XU`�MS.�6jP�9`��TDT��G`~�A>�j� "��'��4$ZO@N�G�"G�U����ePp��e�CN>�G��l�l�iGGROU�W�ª�S� >�MN�kSu�eSu�e`SpW|g|�i�cHR.RpG��z��0CYCc���s�w�cȱ���zDEf'�_D�^�RO�a@s��q[f���vV�Oı 7�%�6��tx�?R�uf��F��m� /k��N1��6�O0'�mB[� PER9�9T��l ,2����5��fGN1LhR1k3 
�-NO��/Am٢��m�����P����CĠ��������O0�nH *�LMm��$U��V ��<A�Z��Ǒ�@N�������7|��8|�9|��~���1���1��1��1��1�ɚ1֚1�1�2R��2����2��2��U2��2ɚ2֚2�U2�3��3��3�����3��3��3ɚ3*֚3�3�4��J!�-f��ao � �$f��VIN�VP�LCWAR�CWqS�T����R��+�FA�C*�SE��$P
 1
�2�������8�<B8��EXT�Ѣap�2��F����U�0tǍe��FD�R��qTZ V�Ec�D1��XR�R�E�F��/�OVM�C��A��TROVf��DT� �MX��ʰ��[� ���IND��
K�5 �0G�z1��
�� #�	�D_��DRIV`�b/�oGEAR�AIO ��K��N�0��EF�F��:`�a/�Z_�MCM � �F��URbr̀��!�? Z�p?(��@K�EE %��Q�!�P��sO���P~]q$VARI��>�X�UP2�t ��#TDPE"}�Gp�5���1_Ti�B;AC�2u Tb�"��4)�:%`cB����IFI��- M�h�����P氯`�aF�LUIWv �8�:P URS�c`���B�1XP} J�EMPd�p�"$Y��?xe�qJނ073VRTU��@x$SHOZ�L��ASShPB1�P��BG_������񢓻񯓻�FO�RC�F�dw��FU�1�22�BR��,P�x |n[�NAV�a�Y�ʉ����S��c$�VISI�пSC�R4SEC��?0؂V�O�$����R����$��I��۰��FMR2��y ��:`�r�� @��ǽ�������������_@���LI�MI ��$dC_L�Mv֛߭�DGCL�FV�|�DY�LD�5�y�5��p߂�>�M�Z`KbzJ $� ��S0�{ P�c� "C��$EX_ !( !1n0�P�aj !39+59&�GtQΤ�| �[�bSW�%ON� �EBU1G��!��GRGpU@mU�SBK.qO1Q�7 :�PO�)P� �Px%� M��O]t֤�SME۱����=��`_E �} ��P��T�ERM	5~5�O�RI�105�QS%MjpO��0�5f���`Q8�+6 �U�PC� �� -<��b}Y� 3�0�~�G�:�ELT�O.��pS(�ONFIwc�1��!ް74�4�$UFR���$��1�0e?OT�G�PT9q��CNS]T�pPAT/Q.DOPTHJmq`Eƀ8�q�r�1ART`�5p�`(B�2RELrJ�qSHFT!R�16A�dH_��R `cO6 Z0$i7�@�_� ��H�s�q�@I�@\U�R} ұAYLOACDYN_�F���6A8+��PERV��Q O�HU�G�prBL����\U����RCE��ASYMFLTR�F�1WJ�7U�Q�EU�`A�YO� aU�T�pQpdE�PVzEPSP�S��Q�GOR�pM�T` �!�ă�"�&�5@�0�q# H��#�� �B�� `O�C�1�!��$�OP��!�c��X����bRE�`R�3��qf�Ѳ7Be?�R�4E�e�h|A��e$P�WR��d�l4PR_`ycYD[ jt�3UDU⸰ Na�2 �y��$H��!CpADDR��H�!G8B\qQq�Jq��Rv��� Hc�SSCv���u����u���u���wO�H�SCD_MN�� q`����`#QHOL������f�� ACRO* �1>�ND_C�s�0Qt>`GROUP=#Bb!_*�;� Ca1{��� _���i�L�i���j��� i���i�����At ��>M"SAVEDd�փ�t�T�s&c� $P�q`_DZ�� ���r/PRM_;Q�&a�PR� �� � �?�D_F�$$CL�S���3`L�^L�_l� O�_ZN�_Zeq��2RdC�@UN�TABC��J�����0V�=1S��ʖ@�$S�VGDLY�HS�SGx$�p�� 񨻰t)*� 3�� SAG� �{#AH�L�0S_cR��_rRlO���_Rƙ_Rә_R���@/�����/5_HTTP_1�H��w� (�OBJ� lJr��$��LE'C��p����� � (e�H�g�_L�T�#�qS��C)�KRL�i?HITCOU���!x�L��`���U���`��`SSP�δJ_QUERY>�A���P_WEBSOC�z�HW��2)a���p�PINCPUM"[Oƶ�Œ۴�t�ޱ�tޱ�� �IA�_CHKCM]� �d�0�PvC3��ܦ�R����NTL�pr`_R_Na;   :�N�N!�0��R2ȮQ_��tV |�S�A6��IDw�VA.�{��pDI��UMMY4;���áƹð�I�PR��U����r|q_� ��������dQ֡őS�����=�6�O�P� �����$I�N��E���"��OT�H	pN�A$WA�T��AF2���$�B������,�S_WCT_�0S����Ik0I70T/�P� �� ����R�R_BIC'�BYP��` �q3�8	p&`/�BT1��`�BT2X�5@'�D �	��"� , s$LBd/ 
$F��5 �㓃
Ja��3� � 8�p�0���X�B��MATRI�XT���BL�`Qr	�Fq 0�� d ���) K����UvSHA1�IZk����$LNT��CH��V�� 8�sq�Ǡ�� <�p� ���0bF��CPDN�! Ap`iT�X����1G� 0`���6T	��� D���(�:�rL��	�ROB
��� ��p!/A�����SL�:���CAkLI��DO �IQK�~�3PO�S�q�  ����BAO@M��0Ǡ�	��0��q�.`��$BI�A�1�QQ	�l�N~^@H � L�p�`i��U��PİICFIX�0E��#4�r8J1
����4�АS�P �1����3���Au��0_HA�N�P� �P| u�x`S��3����1uɘ�Z�X�T;POA<� SKURAN�3�q$RE��H]P2�S��% 9��ʂ��,�O���#)'UBPR�1��/ � k�-"�d%��BO�W�� X��p3љ����LSc��� _a#%�M��k��s$� LIC 'p7!Q�2�eEh��&qP���`�&OSG�>YSWARB��QEXZ�9����75�CH_@NRG�`LI<0�V6ESYN,�TEgSR_@�u7H_���t8ESѱ�CX��Rf�<IDf��5UN��X�%SQ1�=�&�@�0FC�NOK� �Of��7�HR*CR~��_G��L? �u����SFp|Q6`A�er�4�"|? ��� %�7�L�� ��C'�@���pARGIB�L_�N���=�f�8ħGR �GP�yq�F���J�B`Vu�K��H�LAj�h�xU�l ��A����  �~�O�T���r���F�U�RaPˡ�U��M���XU*�@ � x�Nb��8�
��%e}���7�϶���8���e��<Ǡ�����KA ���0�REA�tC�Ѻf�1]� )0ApqHwR����ST%b��dt����R�� =8�U���� ��R	ML���X���Ss��ECK�sgOR�B�԰��܁+��_T� X�3��P}�%b;3��PREFQ ��J�p2�_�  ���P���d] or҂i�ETHO��!"PL�#A��O<BW��SFI=OwPTENC/��WT�]�K�БU�$C�;2�БVUW�TPb�� '�@�TF��">�2$&˱MY��S#�� ބ�avE�C��B�O����DU��O:�boMY30~���ٓ�3��J����E���3����6իҥ�5������	W�T�6��	�Ė	����P҂�Wd�E� s�J�$$��_�Md_�vb(�#�]�����Pj�^��ȇ�zBC3D�_�$����xTP�GL�@AD���I;NI#VOX��ou�֠AZy]�0 ����z����1K�OB2K�1_SP1�k�2p�3p��2m���~�����R�PT�ĵ��Ϸ~� ϳ��˷�ٶ��W��_�Y�EXTRA1$�r/�2a��pRY��q8I���� �Xy|�"�J? APPEh��S@T��FL���w�ZZ����PA���MEMi��=!���R%���]��ZEpf�_�����h������@�="���`Z(����tR�����b!���]� ��C8���6�Y!�Y#n0SIV��E 2p^  _���s���u6�^�����`�&�����]�� ?p�� b#֕�U<��<0VERT� ʃ�q�$0K�	�LEN�����A��Z��MG@��������b Xy����Y��Z�rTOT &�������p� ��!��q��,r.�L�� 4��N�8�A��`�Rp����r�� CDPe�?�t $���Xx}��ERG�P�Ā��n@��[r��R$��Z�D��UE3p��.`&��!�GS����Y��Y��YIN���m���N_X�Y#!I�q�Z�G ���m��]y��V�P������հ��p�[)$ANALY|�@�2!�r� ��ձ���,Ӡ����[��[pnx� �  m� ��� ���}�� �!���I��BGD|F�� � d �aMP�$FI���-;��RLSF?0��"�5TA}I��BUFEX�Qp��^�&"�A� |q�l8&��ME�t��PmI�'SV�(SV�(�CO�)O�(PAT��`).�b�:�b��s @$!ۥ� ��P&1�XDZ q���z{kDn2$TE�q �Qh;���s2y4FLr1�!N��ŀlpT��u��@�'�@���U�P��E۠�b�`VR�WRT�7LNTK��7ARCTOOL�ۡ��A_I#"_C�Zn_ � ` $Z9�}��dFA:��5 TOK�0t1 ^@��8�TAeDnfC.RVE3�D2�`'0b�$�k��D�CPAH��s2
$F�E�0pO7LNK�P���p��0Nb�Pa��; _�2Q7$UP� R���@SLAVE�A� ��O9T4T1WTR,r�O_+!ASޡ� TC@L\�
�N�q3$���pRT�p4��C�p�C��H^/��Q��S��O_U�ܣ�AB�Q.��a�U�`�V�QTRTP^��b�U��a�V&bf'.z� �� XC@IPA9D�Wc_NE�A LAGx�Lp�P-�vf����qF0#�$FO�CUS�@�p  �ITEM_AC5�O� liEŀM`�L����eN�acFpP�dELAہ�d� �F'�$Hc�uR�EPu��ar �	���j�d�dP4��Wu�`Uu�IRCA�D�i�� � T����IT�C�A�S��qC�p�|�Pv��vI�DG8���DAY_pxNT��r�w'R87�r�wSCA�p�w�CLEAR�q����r���a�;\t��hu~r�N_PERC��tp�r�q�`��i�] ��1`J�q'�_OyF�x��2� $0h-qX��a�zP$ކ���`LAB ����`�U	��`�b���կb�U.BRZ��T� H���CURR_UR�!��$AL+�N9U�Q�ISI���Ώ�T_U�s��KY|�B8 ���J�p�a�S`$��F��R�pR�U��_|0N�Pȋ�2QʑJ�2֑FL����p�C둷��1�UsJRb�uQ� ��pF�1�0LC��G���J7b�>�$J8�@�7_A� F�[�7��<�8r�?�APH�I��QJ���DS�B_J7J8A4B�L_KE��[@��KARELM^q k�9XE�ONR;WA��_VA����$N�E��X�y\�Ģ�J��cҪ�V��&�C�T^�0�pe��LD�*4� x��P$�N�TDN�G�E��OR��Ô�NTMO��T�lPD_�: S�PR�OJ��TO������LGK��ȋ $�yL�а38�V���MR��sP��FD��I��������Pp�`� ��MOD�� z��z�sPz�#�z�_��z���~#@RO�0MB���0����Fy������4(�C!
� �0E����sP�#�$�I�.����_�0�T"��R�P0 �cZI���c�aLN4�j
��A@pDE�9RD0��i�I����@L�����DAU��EAaD��
%����GH"ܿPBOO�A��� C�RL`IT0�30�P�VRE�`G�GSCR �ȳ�QD�8�0'�U RGI:Q] �{�V�S���|$QS���TW��Q�ԊSJ{GM��MNCH�D&NFN����K�x���UF��0�FW�D�HLG�STP��V����7��RS�HELc��0�V	C�]�E�dN�����UF!������:���S�G��SETPOb�r�]�����av�EX�WTUI�IS����pS�����@� �-� 'Q�	 d�!d�N���#Z�Q�ǴAV� =4;��D�CSB�3i3O�O(S�sF3S?��IGN�'P>#p�1��DEV���LLy�ֱ��r�`�4�>qT�$�5��r�>4sq]�A}` ��k@�@^a��]`�y`S1%2%3�!ځK�`� ��y	"Ŵ	UF�
Tu��a�ROSpG�[�z&+ST�PR��Y���!� �$p0�$C�+4�FF�'�&��K�a� L_z��X {f�4|`za��N��.4����c�_ � � �0JE�KC ��MC��� ���pCLDP�Pw�TRQLI&����9~4�FL��}1��3;�D��7R�D�5�4�5ORG�����2�ȊO��D�E3�Ao3�� �_��4���4�5&k�PT�0�B	�1kD}sFRCLMC�DHO#O�I4qCP�M���nQvP�ѠͳMAPi��p҃��U��T� ��E\�ja�M�FRQJ�� �� �yHRS_R%U�&1��A�p���FREQ��9�$<� a�OVER�`��q`H&�P�EFIp%1��ϵn0Q�>D� \�QQ[�s$UN ��?_�&�PS\`Ր	\S����D�b�S�CU_p�A�?( 	�4��MISC�� d,��N!RQӒ	�`����pӐEf��RhAX�w���UgnlEXCE�Sm��(bM��0a��>�9bw��(bSC�O  �S���Id_�ՀCh�p�klo~hn0KbK���Rb��FB_$��FLIC4BQ�Q�UIRE���9{O�H{�W�ML(0MJ�� V0?�pK�Da��Bۀ�p�D�"��$T�1+���<A�CKED�qh�c$c�6�tINp"��Y _�  �� ��q9��q)��7���h.�N�C��n0ND�фt�1`ݻҲ�)���D|����INAUTt� ��°5���kN��z����q�t�PSTL�0a� 4א�pQ&R�I� Q%EX	�ANqGƲ�Q�QODA!V��5`$ʠ���MFF�*ŃVw)'2� 158t����FSUP:66@�FX͐IGGC� � �_�'3z�ȳ '3��'4�R�"���  ̘� ۖ�`8�A��QCTI��@�a��M��n�B� t9�MD9�I�)G�WR��AO�qH���R�DIA� R�ANSW��`���kR�D�)�AOR��rk�1`� �`C�U�V��c@%���_�@0a� �? Y#F�L�@в�.��P�h��
�P�KE��;$�-$B����Nx�ND2�BTAR��2_TX04XTR�AW��B��pLOD��1`�b���b������ʢ���� ��M�RR2,e� �0����ApA d�$CALIK`��G�
�2Ȭ@ �
 RIN
���<;$R��SW0�DA��CABCM�D_Jpe�?q�PF�_J3l�
f�1SPYp8 �P	Pfč�3��ϡ� �P���J�C��2BhAO�I&�aCSKP �:������J�b�Q��,��,�"��_cAZoB��^�EL�<�§AOCMP �a��Q��RT	Q�ӧ�11�����q 1�ػ :��Z��SMG��*�v�DJGN0SCL�`��SPH_K`���T@�P��RTEIR@���� #�_	
]1b�A���#b<�sDIt���23U��kDFװ]�LWc�7VEL�1IN/2� ��_BLW�R��'��HA~����MECyH��DTSA_@��װ�bIN�QQ1`�ʢ��p�Q@��� _` ����D�q����b�"�T� ��DH�`��0a��$V�����ӻ$���gQBRD�$TA��R��1`�H ��$BE�p�x�_ACCE��	����A���IRC_=��tO�NT�Q{#$PS�`�2Lװ��s ����B���J���;D��;3
ې�a_!���l rbU�P��_M�GASDD�=�BRFWs0+��������DE�PPABN6RO �EE�! ��0"�!�A�`����$USE_���2S]PkPCTR9Y� ���nA J!YN+`A �Y��i�YM�Aա��� O��-�INC�����Rb�'�.SaENC-�L��R���Pd��IN�"I0
�,���NT~��NT23_a�BR#CLOr�BR3 yPI�p �c=&g���`��� ����aC�&MOSI�� r�raSbPERCH  ��wQ"� �' ��#�@"�D�@��|�C
�q ��A
�%L9���g��%��8@*;6V&TRK �QAY���#�ak1
z5�o3����a�PMOM��Rb�b@Ϡ�d����3]۰DU�&�gS_BCKLSH_C
�5�@{& xPa�SC�&Jp$�CLALM$Q�0A�XECHK���]�GLRTY��D�����q*�_i�p$_U	M�C�FC�C����CnEPLMT��_L��w��D�q�GE�MP�K �@���E����Au0LCT�(PC�!�(H��8fp��ECMC��� .�CN_�N���V&��SF���)VC�����wQ
�U{XCAT�NSHi�¡� �q�1������А 3PA�D�_P�E�3_����r6� ���3�d�EJGM�T1A���p|�W(�TORQU5 ��n#�9� )r�")�� �b_W�5k4�ѐ�tP��u��uI{I-{I��F3�
q��lx��� VC��0&�4�s�1�~� �љvJRaK�|�r�vàDB���M��àM��_DL��2GRVt�������qH_���s> �E�COSR���R�LN�pu��u|���w���@w�Iq����gq�uZp��&�qMY~��^�L�|f��THET0F%NK23��<�{��[CBA�CB{�C�AS�f�Itt���t��A�SB��L�GT	S�C��na��]cx��Ț��$DU�@@7�"�����Q�!Y_WS�NE3�*AK�D��B�_�0�A4��]�f�D�O�O�LPHR�;�%;�S�u���� ����;���أª߆]�EV�Vt�q�V��UV��V��VϫVݫV�V��H�����P��a����H��HϫUHݫH�H��Op��O�O*ɕ�O��O���O��OϫOݫO
�O߆F;�a��ɡ����r�SPBALA�NCE_���LE6��H_4�SP�ᒆ�ҡ�Ұ�PFUL�C�@�(�@Ұ��1=��UTO_}@�E�T1T2����2N dAV ���ѥ1B� �(���1T,0OV���>pINSEGV_!�REV��_ �DI�FW%'�1��T�1�0`OB�HA!��7�2�` oA �LCHgWAR�HABda�5��_ ��A���CXx1P&T��V�b�vЇ� 
���a���ROB� CR2��R_	 �C��_�b�T � x ?$WEIGHu�#$p��`Iu; sIF-� LAGf�ERSf��fBIL�L�OD�0b *�STD��*�P��H@+� ��(`�����
���<g�a  2�m$/�/DEBU;�L3 {�=�MMY9����qNNc���$D3Ʒ!$��`#�   �DO_��A�� <����H�AgS�Be�]�N#�8_D g��OU@ ��� %�@T����AT����TgICK<�P�T1 %��0� N� p�,� R@g`�`�� PROMPuE~R� $IR�`�e�@�0.MAI��p�1w_F����1�@R�CO�D��FUm8�ID�_� J�����G_�SUFFIp h@�\�DO�0�Ь_�GRF�`� ���`�`�a������H6�_�FI��9�OR�De� 	���36�*R�e $ZD�TQ	����4 *�L_NA�A� X"�DEF_Ih(X"�t$�l��v���#��%�IS�$��P$0��#��r$�Q��4�Q=Rv�DPt��24��D�`O��>#LOCKENa������!��UM �X"��#��%��" ��3��#��$�t� �6�!�k��a�X"�@�#��7.E�[ P4� �$k �!9���Wi8hE�_3��TESA��( @�LOM�B_�B�G0*�VI]S�ITY*�A�a}Of�A_FRIqӌ�C5�SI�!�A%�R�� �G� �G3��*�WB�HW�K��F�p_9Y�EAS2��a�DP3`/0�F4�I5�I�63�ORMULA�_INaaTTHR.2���GH'��:����8��COEFF�_Oz���Tz��Gd&a2�S;���CABЄ��$dS1�����G�R$� � � �$_0��-Xj TMR7jd_5�g3�l6�ER �TH4G$���  j�LL�'0SR�_SV"4�h�P�E�����T��� �\bSETU�#MEA� g�p+������ � <`�� ��PCq��Cq71Nv"]"� 71S144$bAQ�~s�00�!�/0�{�7�"RE�C!HqDA�M�SK_��Pd� P~�1_USER������t����p��VE�L�r�p����u`�I<1 ���$$C� F����5���&�� *�RS�B4��@�1N��$AAVM{@K �2 5�w �@�5<�䊏������ ���	܀͍����6��ޏ�� �̌?�K��ہQ���������7 ���ɏۏ���@�'� 5�g�u�k�����Юd��B��P` 1S��? <��� '�9�K�]�o������� ��ɿۿ����#�5� G�Y�k�}Ϗϡϳ��� ��������1�C�U� g�yߋߝ߯������� ��	��-�?�Q�c�u� ��������������)��CC_EPL�M��,����  md>�ING��U� =�)0qP'`l���y�o_CRCR0CO)`���.����P?<5��� ٟ ��#LGYk� ���p��y�������UP$cL��  }d�IOCNV�a
J��U�P�pj����ߣIO_# 1.q�P $���6����~6�?��L� �����//1/ C/U/g/y/�/�/�/�/ �/�/�/	??-???Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OqO �O�O�O�O�O�O�O_ _%_7_I_[_m__�_ �_�_�_�_�_�_o!o 3oEoWoio{o�o�o�o �o�o�o�o/A Sew����� ����+�=�O�a� s���������͏ߏ� ��'�9�K�]�o��� ������ɟ۟���� #�5�G�Y�k�}����� ��ůׯ�����1� C�U�g�y��������� ӿ���	��-�?�Q��c�uχ�>�LARM�RECOV ���p�y�ZLMDG� �u�LM_IF j�q�d&PRIO-�230 Ethe�rNet/IP �Adapter �Error (1�) st 2SS�W0H�3H�)  �11�p�x�d  �NTP-213 �App1 BGL�ogic Not� Running� (BGMAIN, 46) U���[12] 85]xx�����, 
�� �����߀�'�$�3,�Scn��i�n�� Mod  �L�G1L� WOR�LD�m�x�$W�AITPATH � 231 3 B�T0^�Z$ �PAGD ��~�($�6�H�e K�[���1�\NGTOL { ��	 A���b�t���PPINFoO �� �����������   ��������6 Z DV�z��������4�(:L ^p����������PPLICATION ?�������SpotToo�l+R�7$ 
V�9.30P/15���
39104�7?"Q*F0w!d/1�31Q�O,F/X"7�DF3L �7#Noyn�P*FRA�� Q����_A�CTIVE��  �#[�  3UT/OMOD&0��Y��5CHGAPON�LH? \3OUP�LED 1��� �0�?�?�?;CUREQ 1	�W  T�9�<�<�	O-E# BD����2^	.! �Wel��ASW��4��	SWTO;PKwFHKY;O�� �?O"O4O�O�O�O_��O�O_$_*_@N�SD�Handl��aTH�5�2wZHT�A��<_N_`_�r_�_�YSD�Dispens�$ODI�%wDLHL�O�_�_o�o�o�o �o�o�o�o�o+ =Oa����� �����'�9�K� ]���������Ïɏۏ ����#�5�G�Y��� }�������şן��� ��1�C�U���y��� ������ӯ���	�� -�?�Q���u������� ��Ͽ����)�;� Mϧ�qσϕϳϹ��� ������%�7�Iߣ� m�ߑ߯ߵ�������0���IC�5TOL�(?�:3DO_CLEA�Ni?4��NM  Q� �?�� ���$�6��>DSPDgRYR��5HIF0��@����������� �� 2DVhz�8MAX ��Gc
52�X��na�2na>2PLUGG�0��n�3  ��RCY�B���������O�b�t�SEGF `0�@@R[���������"ULAP��Lc6/H/Z/l/ ~/�/�/�/�/�/�/�/|?�;TOTAL���6s�USENU
�; AHq?BB�0�RGDISPMM�C�@VACf�@I@t�4O}�j��3_STRING� 1
X;
��MQ0S:
N�otAtPerc�h�6IsItS�af\d�2	CC_�Manual u�p�4Cycle�Inter3@tu�sASel Pisck�8PBDro4D^_GProc�8yE? W Seq#CQA�Cam �R"D�E2��HTip ChaWnge�@l�2}@�ductionS�taJCChut�H�1QAEcho� Op�A VToo��@�B�1Auto3_C�1�6  Q�;�@_R_d_�3I/O SIGNAL�5�Tryout� ModEI�np�PSimul�ated�BOut��\OVERR~|� = 100D�n c>A�8}@g� Abor�S RR�obot iCAl�oWBe isYo�QQOn�@p `/Weld�S�T�E�$BHeartbeatr_p_�o�o�o�o �o�o�o�7���;>��_ITEM�F Yk}����� ����1�C�U�g��y�������1qWOR ^�;فM����%� 7�I�[�m�������� ǟٟ����!�3�E�W�PO�;%A}�� f�����į֯���� �0�B�T�f�x����������ҿ���x�DEV��!����H�Z�l� ~ϐϢϴ��������� � �2�D�V�h�zߌ�>��PALT9}�� �������#�5�G� Y�k�}���������������1���GRI� �;i���C����� ����������!3 EWi{�����W�O0R9}��� 5GYk}��� ����//1/C/�U/g/y/�PREG �޲ %�/�/�/�/? !?3?E?W?i?{?�?�? �?�?�?�?�?OO]��$ARG_ـD ?	���`A��  �	$V	[�tH]tG�W�IS@S�BN_CONFIQG�P`K�A�B�A��ACII_SAVE  T�A�CS@�TCELLSET�UP `J%HOME_IO]~\%MOV_Q-_3_REP~_IJUTOBACKP�`I�A	M�C:\PROG\��' � @ ���Q h�,�@ՠ,`�'�'�� �[�@ �21/05/08� 02:24:16�&�H�-?oQo~o<uo�* ���o�o@�o�o�o�&��o M_q���2� ����%�7��[� m��������@�ُ�����!�3�E�� � �U_�S_\AT�BCKCTL.T�MP TER��.}Tl�RBT01���������Ɵ�_TOE�X�B �^E��� AcCz ; Bi  e�E疿GRP 3`E��@ t�V �'�T0���@�C�Z�R��M`58��z�9�EA��)`A�)d�D�1��Đb6C%M�|=�o� �(.R��P�b�� h��� �f��  ��٥G�#��-�C<��L�^�t� "���������ҫ迷�������PORT �[	 b�Ae�Ts�_É��A��zA`ϾτƊ�������WRK ?���U���C
��CWߖXI�NI��e�F�SMESSAG�@{��A�P�C�A��ODE_ADP�F�E5Դ�O���ߛSPAUS� �!�`K ,,		h�`E�+��K� 5�W�Y�k������������#���Y�������TSK  �P��h���WRCV�_ENB�@�M5�UgPDT��y�d����XWZD��{��J��STAx�`A��RA�XIS�@UNT S2`E�A�@���VEl=�y�s�Q� � ��o��V�� :XF8)q���� `O� �4� P�р� ?��  ������0��n	47� c\_��U9�ݬ�q�ؕ/1ME|� 2�D	T�P��A���A�P�A�e��@��Aٶ߀B}�-:��G:��:��v�9��T:��F�:*^�-=cK�'��/�-L5��&/XSCRDCF�G 1?��P��E�B/3?E?W?i? {?�?�U�?:Bx��G ? �?�?OO%O7O�?[O �?O�O�O�O�O�O@OzO�W�QGR= �����Sk�NAME �	��	�TV_E�Dw�2H�
 ��%-q�EDT-�_�)%�_�_� *@�U�QXR�_$��ϰ�U�_4o� ��"e20+o�_xo�n�_��Y�To�ooo�o<o$c3p�ogoD�o� �[� ��o�oz$c4�3�W㏵�U�@W���F��$c5�� �{m��.��U��#�j�|����$c6[�ˏ�� �����6�H�ޟl�$c7'���t����P�@������8�$c8��@�R��6���� ί�v��$c9��/��S��6��SϚ���B�п$aCR*ob��� �Ϙ����d�v�ߚ��PePNO_DEL�$_6RGE_UNU�SE"_4TIGAL�LOW 1���   (*S�YSTEM*�#�	$SERV_G�R\R�W*x�RE�G��$��]*�NUM�*��]P�MU�о%LA�Y? �,PM�PAL�5^�CYC10�_x�a�e��ULSUW��y�x����L����BOX�ORI	�CUR_����]PMCNV6S���10��?�T4DLI�����Y�	*PROGRA���PG_MIe����ALo��������B����$F�LUI_RESU`}��);MR���P5�5ߗ��� �����!3 EWi{���� ���////A/S/�e/w/�/�/v�LAL_OUT ���c7QWD_ABO�R�0��`Q� ITR_RTN  �D����� NONST�O\P'4 8CE?_RIA_I��'5�p0��Z0FCFG HZpDgM�y1_PA��GPw 1�;�.��O�?�?O�;C��  0MD� D_@ DB@#F@U-J@7B@@F@JJ@V~�D]F@gJ@qB@�zB@�B@��3D;�� �NIF@XB@f�J@t�@�` D���@�� D�F@��� D�B@�  �D�J@��@��@���F?�O�?__T%_ N|2@�2@�2@_�� C�VP�VPU�VP�VP�2@�2@U�2@�2@�2@�VPU�VP�VP�VP�VP�2@�B_T_f_x_�\��HZ0HER�ONFqIG ?�QG_P�;1�; o��� BoTofoxo�o�o�o�o��QKPAUS��1��p3 ���o ���o4DjP� ���������0��T��lM0NF�O 1��>�0 � 	�O������W���4ſ'X�"���²�Q���5#f��@�2��ĐbKC%W(�=��K�\��$��Eټ������D�J�%4�+ɵ���B�����1���H 3�[��f��Fm�f�Z0�O}1�?�8��L_LECT_}2��1�"�7˗ENo�'5���璤�NDEӓ�!ۗ30�12�34567890�;�j2�ѓ29�K�f�
9 I��/  )���� �̅������ɯۯ4� ���#�|�G�Y�k�Ŀ �������׿���T� �1�CϜ�g�yϋ��π������,������2"ۛ ����IO $$��f�&6�������߈�T-R�02%`�(��ف
�f�(�a��`�&��P�y�CO_M�ORm3'�< ����aB���A?G�F�����A@�D �����������;��Y �w�e�����������T�3��(��,e?�A�A�@T K"L��H�#Y1P�*۝��8�O���@�
 ���7� �"�B@�=��=�@� �wsja�PDB ��,�,�cpmi�dbg;�;`�:���}p���/  ���/�����g/��D/mgX/�/|/��f�/�/F��/�u�d1:?G?��`D�EF +>���)�21cW!buf.�txtR?�S?c _�MC��2-gn�df�? d�3��2.�=���E C=B_@��CI�BI����A��As���A�B%��JA�8�B��j��B���B���LB���C��]`Cs/C��tZ��D�?E����D���E�aE��E'F�@��D\}#F<@�4IC���?6��E�Pr�_��H�A��XA_�M�2��0`ܫDu�Y�Y���Y�  @��M��Px�A ��P�U��CD�P�N�UUD�nD�t]E;� Dz�  Enb�N^�8�DD��;;E�` E�@ E�4A\���  >�33| C�I�@�n%��5��I�%AG@�=L��<#ס��4P�o�Χo��d~�S��1�U�1�W�Q�_G��$J��<J\2g=oOh�� Qeeowo�o��o�g�2�RSMOFST �)q:b�p�P_Tm1Y�31`�A�P�I�`�A�MODE ;2۟��Y�q��;��r��w?����<�M>���;:TEST�k1/q>��RՒ3(���#G4�p�@��PU �Q�qC�PB�T�B��CCK�8���Y�:dڡ� �q��Mq������*��I�4�?��Z҅5��Q��1����T�_�PROG ���%	ALTM�ASTER A��r�.��TD f�$��R�INUS+� �U`��I��KEY_TBL S g`�� &��	
��� !"�#$%&'()*�+,-./012�3456789:�;<=>?@AB�C�GHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~�������������������������������������������������������������������������������͓���������������������������������耇��������������������P��LCKR��I�R��STAT����_AUTO_DO ����$ͲINDTo_ENB�� Ͳ�F�׿ɶT2��&6Q�SF��6�����U �(UT1:�E��@��j�M�GROU��7��=�)A�B&��C���B��~A�2`��.7���@�B���b=̀JY��E�� �7 !�Y�9�K�]�o߁ߓ� �߷��9A�p<B������ľP`�C�f�GCP�RW�`��.�;�M� ��m������W�0�����J�TO ������TRL
�LET�E6� ��_CU�RSCRN 48�� ��?�Q�c��u���YT_�EE�N ��k�csc��U��MM�ENU 19g <�l%�o� ��@3C|S e������� 0f=O�s �����/�/ P/'/9/_/�/o/�/�/ �/�/?�/�/?L?#? 5?�?Y?k?�?�?�?�?  O�?�?6OOOlOCO UO{O�O�O�O�O�O�O  _�O	_/_h_?_Q_�_ u_�_�_�_�_�_o�_ oRo)o;o�o_oqo�o��o�o�o�y��_M�ANUAL���Z�CDP�:�e�g�"�+㩇��?|(����EtI�;O�B8�*�?i���re���j�DBCO�RI�G�碹DBG_E7RRL�<�˽�a�O�a�s� �q�NUMLIM6�������DBPXW�ORK 2=���>�ӏ���	����D�BTB_�� >�+�e��e��#qDB_AWAYb�pq��=���q�_AL����o� ��Y �����q�� �2?�}, 
�`�U��+�5�_M�IS��~�@�C�OoNTIM����3�e���
��̗MOTNEND�����RECORD ;2E�� �3�U�G�O����U�S� '�9�K�]���e����� ���Կ�������.� ��R���vψϚϬ�G� ��?���c��*�<�N� ��r��ϖ�ߺ����� ��_���8��\�n� �����%���I��� �"�4���X���Q��� ��������E������� 0���qWi{��� �2��� A,�w�T�� .��d/�=/O/ a/�/�//�/*/�/��/?�/�,o�TOL�ERENC|�B��Œ��L���pCS�S_CNSTCYW 2F���<�?Ò�}?�?�?�?�?�? �?�?OO-O?OUOcO�uO�O�O�O�O�OX4D�EVICE 2Gh; W�_4_F_ X_j_|_�_�_�_�_�_�4�Y3HNDGD 3Hh;��Cz�ZБ�[1LS 2I	] �_Xojo|o�o�o�o�o��_Z2PARAM JR}1U1UFaZ�X4�RBT 3L���8�<&__� 7C�wv�b��q/C�  eu�npW�,V�PvD [x�ks�A��E��vW�I~�[wmu�L0K1�u�x�qT
sVq��x�wp4�o4�StH[w�wpd��i�X�W���L{a�[w�A�ft��Öu  czVp�f��Џ�� ��ˏݏ��N�%�7����  DV� D�`Dl(�� 	 �B�ffAp � Aə�A�3�3A���BfAf�j��b�Ֆ�tC���̗�#�B>ff�B<�|I0|������şן� �U{� ��� ��33 m�� _aW h��n >s`�r���Z������� ��Я����S�*�<� N�`�r���ѿ����� ޿���&�8υ�\� nϻ��Ϩ�������� �>�)�b�M߆ߘ�s� �ϳ��߷�������� �#�5�G��k�}��� �����������H�� 1�~�U�g��������� ��w� 0VAz e����߯���� ���R);�_ q����/�� <//%/7/I/[/m/�/ �/�/�/�/�/�/8?� \?G?�?k?�?�?�?�? �?�?�??FO?/O AOSOeOwO�O�O�O�O �O�O�O__+_x_O_ a_�_�_�_�_�_�_�_ ,oooboto�?�o�o �o�o�o�o�o: OCoUo�Yk�� �� ���6��� >�C�U�g�������� ��ӏ���	��h�?� Q�����ԟ����� ��@�+�P�v�Q� ����������˯ݯ� ��%�r�I�[���� ������ǿٿ&���� \�3�E�W�i�{ύ��� U�������4��X�C� |�gߠ߲ߍ����ϣ� ����0���f�=�O� a�s��������� ����'�9�K���o� ������������: %^I[��������$DCSS�_SLAVE �M������
_4D � !AR_M�ENU N  ����hz�������\a�/:S�HOW 3O � �N/��[ m//�/�/�/�/�/� �/??��D/>?h/e? w?�?�?�?�?�/�?�? O.?(OR?OOaOsO�O �O�O�?�O�O�OO_ <O9_K_]_o_�_�_�O �_�_�__�_&_#o5o GoYoko}o�_�o�o�o �_�oo1CU g�o����o��o �	��-�?�Q�x� ���������� �)�;�M�t�q����� ȏΏ˟ݟ���%� 7�^�[�m�������N� ǯٯ����!�H�E� W�i���������ÿտ ����2�/�A�S�z� tϞ��ϭϿ������� ��+�=�d�^߈υ� �ߩ߻�������� '�N�H�r�o���� �����������8�2� \�Y�k�}��������� ������"�F�CU gy����>��~.CFG P,�6�dM�C:\$ L%04�d.CSV�3 c�="�!A jCHrz���
6������<�7 s�y���$3 3 �R�C_OUT Q�& m �o q s�_F�SI ?L) +��/�/ �/�/�/�/�/!??.? @?i?d?v?�?�?�?�? �?�?�?OOAO<ONO `O�O�O�O�O�O�O�O �O__&_8_a_\_n_ �_�_�_�_�_�_�_�_ o9o4oFoXo�o|o�o �o�o�o�o�o 0YTfx��� �����1�,�>� P�y�t���������Ώ ��	���(�Q�L�^� p����������ܟ�  �)�$�6�H�q�l�~� ������Ưد����  �I�D�V�h������� ��ٿԿ���!��.� @�i�d�vψϱϬϾ� ��������A�<�N� `߉߄ߖߨ������� ����&�8�a�\�n� ������������� �9�4�F�X���|��� ���������� 0YTfx��� ����1,> Pyt����� �	///(/Q/L/^/ p/�/�/�/�/�/�/�/  ?)?$?6?H?q?l?~? �?�?�?�?�?O�?O  OIODOVOhO�O�O�O �O�O�O�O�O!__._ @_i_d_v_�_�_�_�_ �_�_�_ooAo<oNo `o�o�o�o�o�o�o�o �o&8a\n �������� �9�4�F�X���|��� ��ɏď֏���� 0�Y�T�f�x������� �������1�,�>� P�y�t���������ί �	���(�Q�L�^� p����������ܿ���$DCS_C_�FSO ?����� P ���7�`� [�m�Ϩϣϵ����� �����8�3�E�W߀� {ߍߟ���������� ��/�X�S�e�w�� �����������0� +�=�O�x�s������� ������'P K]o����� ���(#5Gp k}����� / �//H/C/U/g/�/ �/�/�/�/�/�/�/ ?�?-???h?c?u? �C/_RPI�)ϋ? �?�?�?�?��?	OROX{OvO�SL�?@GO �O�O�O�O__C_>_ P_b_�_�_�_�_�_�_ �_�_oo(o:oco^o po�o�o�o�o�o�o�o  ;6HZ�~ ��������  �2�[�V�h�z����� ������
�3�.� @�R�{�v�����ß�� П����*�S�N� `�r������O4O�O�� ���&�8�a�\�n� ��������ȿ���� �9�4�F�Xρ�|ώ� ������������� 0�Y�T�f�xߡߜ߮� ���������1�,�>� P�y�t�������� ��	���(�Q�L�^� p���������������  )$6Hql~���!LNOCO�DE R8E��"KPRE_?CHK T8K� �A � �< �� 8E@R8E 	 <4��أ t����/�� </N/(/r/�/^/�/�/ �/�/�/?�/&?8?? \?n?dV?�?�?P?�? �?�?�?"O�?OXOjO DO�O�OzO�O�O�O�O __�OB_T_._`_�_ �?�?�_�_l_�_o�_ �_>oPo*oto�o`o�o �o�o�o�o�o(: FpJ\��� ���_�$�6��Z� l�F�����|���؏� ď� ���D�V�0�B� ����x�ԟ����
�  ��@�R��v���b� ������������*� <��H�r�L�^����� ��޿�ʿ��&��.� \�n��zϤ�~ϐ��� �����"���.�X�2� Dߎߠ�z����߰��� �����B�T�.�x�� D�r����������� ,�>��*�t���`��� ������������(: ^pJ���� ���$�0Z 4F��|��� �/��D/V/0/z/ �/f/�/�/���/
? �/?@??,?v?�?b? �?�?�?�?�?�?�?*O <OO`OrOLO~O�O�O �O�O�O�O_&_�/_ \_n_H_�_�_~_�_�_ �_�_o"o�_FoXo2o |o�ohozo�o�o�o�o �o0B8_*x� $������� ,�>��b�t�N����� �������̏�(�� 4�^�Tf����@��� ܟ��ȟ�$���H�Z� 4�f���j�|�Ưد�� �����D��0�z� ��f���¿|�����
� �.�@��d�v�P�b� �ϾϘ��������*� ��`�r�Lߖߨ߂� ����Կ���&���J� \�6�h��l�~����� ��������F� �2� |���h����������� ���0B��NxR d������ ,btN�� �����/(// L/^/F/�/�/�/�/ �/�/ ??�/�/H?Z? 4?~?�?j?�?�?�?�? �?O�?2ODOOhOzO p/bO�O�O\O�O�O�O _.___d_v_P_�_ �_�_�_�_�_�_o*o oNo`o:olo�o�O�O �o�oxo�o�o J \6��l��� ����4�F� �R� |�V�h���ď����� �o�0�B��f�x�R� �����������П� ,��P�b�<�N����� ��ί௺������ L�^�������n���ʿ ���� ���6�H�"� T�~�X�jϴ��Ϡ��� �����2�(�:�h�z� ߆߰ߊߜ������� �.��:�d�>�P�� ������������� �N�`�:�����P�~� ��������8J $6��l��� ����4F j |V������� �/0/
/</f/@/R/ �/�/�/�/�/�/�/? �/?P?b?<?�?�?r? �?�?��OO�?"O LO&O8O�O�OnO�O�O �O�O _�O�O6_H_"_ l_~_X_�_�_�_�_�_��_���$DCS_SGN U�5�(`���`w�16-JUL-�21 06:07�   -d55f5:�1Aa[`[`G � R��:ib�s	"qaeb��}i�ea-a�ul�s������k�o��kcVERSIO�N  jV?4.2.14[b�c�`EFLOGIC� 1V�5?�  	�P�e��0y�0~�bPR�OG_ENB  ��d�cIp4sUL�SE  uLu��b_ACCLIM^_v�Ns�ssWRSTJNT_wv(a�dEMO=|�HqPq�b�pINIT� W�j�:�vO�PT_SL ?	��6�r
 	Rg575�c�74#��6$�7$�50H�1�H�2$�xr��g�T/O  ��h����lV�pDEX_wd�(b[`߃PATH� A jA\ �ASKROUTF�IX\  D_2�1_7_31_0�1_36\ 1�2�7\ 3_03_�24&�ЏHCP_�CLNTID ?<�f�c x�e�}��bIAG_GR�P 2\�5? �'��0�F?h F��.ΒE�֓u��Ȑ�B�  ��B�����
�C_��C��$�G�L*=C�M�JB��f373 6789012345n���w�0� �=�qB��(�B���B��B� {A��HA��33A��A�؏J���[a@�  AB`Ap̡͠��KA�����B`B�i�\c�e�[a
��1�33B,z�B'���"��p�B��B�\Bo��B9� ��� �2į֯��:���>�}5�Q�B��}!��HB1��(�A�Y��G�A�{C�U�g��y����A�
=A��尲��A�p��A�尢=qAߜffA�I���
A��Ͽ����)�ĥ��=���A���A�I���Q�A����U�����=q[�m�ϑ���)����L�ͅ�A�\)A�5���z�A��A���A�ɰ��� ������/�� o�� �>���,�� �J�t� R���4�F�����@��(�:���F��3���,���C���\��=m{�h��>#�
����8b0��7Z�����@ʏ\h����f`@�Ah�Е�����<��/4�9X<��=�+=0 ��;���W�a��_`��>�v�C�  �<(�U[` p4r��М����V��A@[b���� X� ��c�AP[b�	 ���[`Zbg��c�Y�k�g�o��m�?wG+�Y����㝽�G�%�B�\%��9�8%�D$����`%k%3���C�%�"L?(�CM�)W�Ǒ��/�,���/㝏�� ?N.E�  E�lِ,1@22D�?�	`?[a�U?����4[q;�E�:3t!0�:��oλʌ���7�0�D�2��Đ`�C%Nl [`�e��N?�?J?�?�)�OB�9�9=��)���!v��?`O�?�OoO�O�O�O�O퓾�L���#�������P�;����ŕn��O0_�O T_?_x_c_�_�_�_�_e�s�s����_ o2n oUogo���¢��o ��o�o�o[��o'9 Io�oU�� ����#��G�Y� 7�}����c�u�׏� Ǐ�����A�g�E� w���'�9������՟ �-���=��u���e� ����G�᯿_��_,� �P�;�t��� _��������qj��D� ,��-�]ϣmϓϥ� ;����u������5� G��n�ɿ��}ߢ��� ���������4��X� C�U��y�����i? �h��)���M�8�q� \������������������7"[�F=+�ߎbO�Yߢ��$�DICT_CON�FIG ]'����V`�eg���ST�BF_TTS  ���
���VERa�� MAURST � �5MSW_�CF� ^���0�OCVIE�W"_b�A���;UD1:\DC�S_BUY_OF�1_00\PR�OCEDURE �TO RUN TWHE � � �.PDF��/.���8/J/\/n/�/�/ !/�/�/�/�/�/?�/ 4?F?X?j?|?�??/? �?�?�?�?OO�?BO TOfOxO�O�O+O�O�O �O�O__�O�OP_b_ t_�_�_�_9_�_�_�_�oo(o�RC[	`'�/!�_qn_o�o��o�o�o�o�o QS�BL_FAULT� aRj��uLTTBL 1b&{
 (
z��\ n������� %��"�4�F��j������Ǐ��tGPMS�K-w� TDIA�N`c�	n'��'� 6789012345;��/�R�P�w����� ����џ�����+� =�O�a�s�������+��@
f�߯�TR'ECP�&�
4�&� M�_�\�n��������� ȿڿ����"�4�F� X�j�|ϣ���ǯ��9m�UMP_OPTIcON&~��TR[t*y�PME~��Y_TEMP?È�3B�(Y�s�AV�C�UNI@�Y��YN_BR�K d�xEDITOR����2ߧ��_��ENT 1e�Ri  ,&�WAITPATH�  231 3 �BT01��� &;	S?�SSW�����-�]&STYL�E?� S �Y�&�TIPDRESsS_K�|&Tq�?THOM Ev�|������_POUN�C����&CAP_CHANG��>	�&CC��w��0R��d&M�OV_��E&�e&�	�4  020XX����AU��R�����
_ALTMA�ST"����WR_7UPD��B1����#SE��W��=0L)�MPR��|�R MV2PT���TOOLDA'TAU��n�r�{ETv�2_1 V��tEMGDI_�STAl��Y� �� ��NC_I?NFO 1f�۹������`���x`1g�� �P����.
.d�� G/Y/k/}/�/�/�/�/ �/�/�/??1?C?U? g?y?�?�?�?�?��? �?�?OI4!OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_$J�?�_�_�_ o+O5oGoYoko}o�o �o�o�o�o�o�o 1CUgy��� �_���	�#o-�?� Q�c�u���������Ϗ ����)�;�M�_� q����������ݟ� ���7�I�[�m�� ������ǯٯ���� !�3�E�W�i�{����� ��˟տ�����%�/� A�S�e�wωϛϭϿ� ��������+�=�O� a�s߅ߗ߱�ÿ���� ����'�9�K�]�o� ������������� �#�5�G�Y�k�}��� ������������� 1CUgy��� ����	-? Qcu������ ���)/;/M/_/ q/�/�/�/�/�/�/�/ ??%?7?I?[?m?? �?��?�?�?�?// !O3OEOWOiO{O�O�O �O�O�O�O�O__/_ A_S_e_w_�_�?�?�_ �_�_�_Oo+o=oOo aoso�o�o�o�o�o�o �o'9K]o ��_�_����o �#�5�G�Y�k�}��� ����ŏ׏����� 1�C�U�g�y������ ��ӟ��	��-�?� Q�c�u���������ϯ ����)�;�M�_� q���������˿ݿ�� ��%�7�I�[�m�� �ϣϵ���������� !�3�E�W�i�{ߕ��� �����ߋ����/� A�S�e�w����� ��������+�=�O� a�s��ߟߩ������� ��'9K]o �������� #5GYk}�� �������// 1/C/U/g/y/�/�/�/ �/�/�/�/	??-??? Q?c?u?��?�?�?�? ��?OO)O;OMO_O qO�O�O�O�O�O�O�O __%_7_I_[_m_�? y_�_�_�_�?�?�_o !o3oEoWoio{o�o�o �o�o�o�o�o/ ASe_�_��� ��_���+�=�O� a�s���������͏ߏ ���'�9�K�]�� �������ɟ���� �#�5�G�Y�k�}��� ����ůׯ����� 1�C�U�g��������� ��۟���	��-�?� Q�c�uχϙϫϽ��� ������)�;�M�_� y�gߕߧ߹�ӿ���� ��%�7�I�[�m�� ������������� !�3�E�W�q߃ߍ��� ��g�������/ ASew���� ���+=O i�{�������� �//'/9/K/]/o/ �/�/�/�/�/�/�/�/ ?#?5?G?Y?s}?�? �?�?��?�?�?OO 1OCOUOgOyO�O�O�O �O�O�O�O	__-_?_ Q_k?u_�_�_�_�?�_ �_�_oo)o;oMo_o qo�o�o�o�o�o�o�o %7Ic_U ���_�_���� !�3�E�W�i�{����� ��ÏՏ�����/� A�[mw�������� џ�����+�=�O� a�s���������ͯ߯ ���'�9���e�o� ��������ɿۿ��� �#�5�G�Y�k�}Ϗ� �ϳ����������� 1�C�]�g�yߋߝ߷� ��������	��-�?� Q�c�u������� ������)�;�U�C� q������ߥ������� %7I[m ��������!3M� �$EN�ETMODE 1�h��� W ]�]�}�X�}��\OAT�CFG i������C���DATA 2�ji��z*�*�/+/=/O/"^+d^/+��W��/ �/�/�/�/�/??�/ �/O?a?s?�?�?�?#? �?G?�?OO'O9OKO �?�?�O�O�O�O�O�O �OgOyO#_5_G_Y_k_ }_�O�__�_�_�_�_ oo�_�_Uogoyo�o�o�o�m\RPOS�T_LOG l�Me
�'9�[RROR_PR�`%i%>o{Jx�TABLE  �i������kR�SEV_NUM �x  ��s��a_AUTO_ENB  ��qJt_NO'� �mi{�  �*�j��j��j��j��+i�������C��FLTR/�A�HI�S�Oaq<�_AL�M 1ni �2Mdj�W�+��C��U�g�y�������_O�UT_PUT 2�o�Md,z,���d_�I�  �ih�|�\T�CP_VER �!i!j��$EX�T�`_REQ�9�:�l�SIZu�g��STK��X�X~i�TOL  Oa{Dz��A g�_BWD��Ϡǆ����DI� p��g� �STEP��#�\=�OP_D�O��ZFACTO�RY_TUN�d�|�DR_GRP �1qid 	��ӿ|İ~�v�9"��0���7k���F ����ĳ��*�İA~g�B���B���B&��BsqA~���/�@C�BA��9dB27�A��i�B�H@7��W�Pȑ����/͢���cª�!A��2+A�7ZB��OaA`d��/���\c����)������z���{��a����0�B�
 J窚�o�MeA��pB��Ƶ�ϛ߭ߘ߼��8�C�  ��`���W�UUU�UU���<��� E��� c�.�P]���Q*.a��Nȗ�l��M�D/�?xy��Q�:�?>���8��/���J���I\ �������oh��$b�+�ٿۿh��2��`�χ� 2������������<)8�B���.1����VY~� SѦ�{���� 1U@ydv� �����//?/<Q/(�����R/���FEATURE �r�u��`��SpotToo�l+ �(ObE�nglish D�ictionar�y�'4D Sta�ndard�.An�alog I/O��/A� e Shi�ft	?uto S�oftware �Update.9m�atic Bac�kup�)\1gro�und Edit�ing�'Came�ra0F?Cel�l<�7nrRnd�Ima3�<ommo�n calib 3UI�3�;sh�1�?��7coA0O<0pa�neCLty0sOelec$0�6nz1��0Monitor�CJns� t Pa�thNntrol Reliab0^CJrner�@gpA��+DHCP�:�Ia�ta Acqui�snC�Iiagno�sX11�Kis�BF�aults ^pe�nse Plug�-i\splay�}1LicNR�Goc�ume�@View��@�Jual Ch�eck Safe�ty�1�&hanced Mirry@�Image�]Ro�b Serv�@q�]T1s@d�J�V�54o`s�@Fr�0�'�xt. DIO �j@fiT?gend��PE�RLR[m3gs�Zir� J` ꠹*F�CTN Menu�Pv�C�gTP I�n�`fac�e�%G�igE�n�es0p �Mask ExcڼPg<gHT�`Pr?oxy Sv�Tvigh-Spe�P�Ski�4uPN`mmunicW0�@Ux�ur�`�`�O1�bc�onn^A2�xnc��P�@ru�"�z�pe�Q�PJU�$KAR�EL Cmd. �Lpu�P�|Runw-Ti;`Env�xԝ`@@+[0sY0S/�W�'qU�R�\q`Bo�ok(Syste�m)�*MACRO�s,Lr/Offs�e`GMH gri�pp�@c�3l�MR�s@oB^Mat.H�� l}1OpSo�e�chStop*qt ^@ڊ�S ;��x�P0�Y0��QSwitc�F1�oBQ.N`%J���׀ma���+pfilď\��g�wo�8Pi Appl��AzA��eE�@p�R��-Tp�}3�)PCM fu	n�w�o T�R�/�d�Ad�r;Q�ri�@qF�g�0Num�P�]A�C��9` Adj�u`p}��� :��ta�tu;\���!Boxp���Y��RDM�Q�ot� scove��!+�eaȐ;`Freq Anlypw'Rem�Nan�'+��7��QrP�Quest��oN` kSNPX� b,��.SN(pCli�O�br$���!2Libr�#�� ��U���oI�t�`ssag���� RZ�(�T�@63��t�GsPr3ed�#z�/I�m{şMILIB��~�P� Firm?2��PκcAcct0|;TPsTX�O|�eln�������  ����or��� Simula(xA�1[�uC�P>Fv�hs0�A]�&��v.?��70ri�P3�USB port �0�iPe`�A��R E�VNT����nexcept�Pl�=���,4hmVC�1rkr���W��@h���y��s�S�ݰSC-ի�SGE����UI�+Web RQ;U���Q� �2p�T�Q�fZDT˒it�*Z�EOAT��`4�&x�����Grid;��iQ���iR_�.��*��Q��r�-900iB/700�~��Gun Ax�`��*� Graphi9c��%DV-�@�BCtrAJrGs~�%�dv�SDCS�@c�k�q�%larm �Cause/j�e}d�(Ascii*q���Load�@�
Upl� &?80\1?0w0cxil�/9kcRe?�62Tgp~0� �*+��c7ere�P C:�+��j���CJl� pAGu`�&����6yc0��n��ЭP�F�os./Gsc�R��Q2,�uCX 2v0a�#�Җ{VmaXPN:a�Q.k�P|�P�Ѻ*�R��Outpul�*A�jtherNet���T�+I�Snifpy�.I��!Ada,�<z@�/ EDA�/�$�Sca�p8ceAx#isNa�A�mm�Q[D��eANUC��@Cr�eRA�@9`��e�A t��p��vte���-�PMC�|�;Paksh�bI�q�/C��o�V�qR R�]�0�Lƃp�en�Q�i�`<��bUtil�H����M���
t���VNR�TJN��OnҀe Hel���H��e㹀b^���o���0�35G�:Y4�FA���Wi�z��asswo����PayId �^"�Y�S�pf����a�^���tr�{+pc�R�pa������W5%�OS �&�eP�j����3ׅ��Z���Av�oi��c�5MqJu#mp�zC��F���_�Easy NoCrml0����Cˀ1 by E-����PEED OUTPU��~��oB��J�s�{nost�^?�64MB D�RAM�O�sFRO@�4�h�b/�}M/yx���allb�@&��R�׀�T�s# ��G%�Q!	
G%k�)k`(MAILE�a'P ����'?"Adp.֍�s;0A?S2��z6�� s���Hig�>p"�6�6ABIC|`��}Inclu� h��?�L�@ar;���0UR��UL �%���OPT���`�&PS�M0p�cro�HW#AY%�g�R�u ����\ޚG���p��Syn.(RSS)G�quiK� �&�7�@������p߽��S&P�e�"texhlVG$�A� d�N�1w%0jo�2
3Te�`��,̨;WTp�e��3
�H4�FTX�S	 dut��U�g�0cap�:˽t�0inf @ͧ�g�c
�dLim *�nS�6�1�v@ K�tes�)�0K1e�F��ldx0	#�{�?� �ϭϿ�������"�� +�=�O�|�s߅߲ߩ� ����������'�9� K�x�o������� ������#�5�G�t� k�}������������� 1Cpgy ������	 -?lcu�� ����///)/ ;/h/_/q/�/�/�/�/ �/�/
???%?7?d? [?m?�?�?�?�?�?�? O�?O!O3O`OWOiO �O�O�O�O�O�O_�O __/_\_S_e_�_�_ �_�_�_�_�_�_oo +oXoOoao�o�o�o�o �o�o�o�o'T K]������ ����#�P�G�Y� ��}�������ŏ�� ����L�C�U���y� ������������	� �H�?�Q�~�u����� ���������D� ;�M�z�q��������� �ݿ���@�7�I� v�m�Ϭϣϵ����� �����<�3�E�r�i� {ߨߟ߱��������� �8�/�A�n�e�w�� ������������4� +�=�j�a�s������� ��������0'9 f]o����� ���,#5bY k������� �(//1/^/U/g/�/ �/�/�/�/�/�/�/$? ?-?Z?Q?c?�?�?�? �?�?�?�?�? OO)O VOMO_O�O�O�O�O�O �O�O�O__%_R_I_ [_�__�_�_�_�_�_ �_oo!oNoEoWo�o {o�o�o�o�o�o�o JAS�w� �������� F�=�O�|�s������� ��͏ߏ���B�9� K�x�o���������ɟ ۟����>�5�G�t��k���  �H590����21^��R782��5���J614��ATU]P֦545֨6���VCAM��CLI�O�RI�UIFz��6��CMSCB���STYL֧28v6�63�NRE6��5�R52�R6�3��SCH�DS�BZ�PLG��LI�C��DOCV޶C�SU6�9q�ORS�R6�8��R869�֧0�EIOM�R�54ɦ���ESET��J7�����MASK��PRX5Yf�7��OC�j��}���ɦj�ը3��J�6Ԩ53%�H��L�CH��OϸJ50n}�MHGM�PSз�MϸMCX�*�m�5���MDSWv״�OP��MPR�����OMAEN֨��0��PCM5�0��j�᦬*���51��5��5�0��PRSa�R5� �J69��FRD��FREQ��MC���S�H93��S�NBA6���SLC.�SHLŷM�窰��SPP!�2��2��HTC�TMI�e�Ơ%�TPAM�T�PTX�EL��5�0%�8ȧƠ��J9�5q�TUT��95��UEVa�UECn��UFR�VC��wVCO�VIPe�wCSC1�CSG����I��WEB�HTT�R6��S�꠶��CGIG��I�PGS:RCe�D]G��H79��H#�R76��8hז ���R85�66�7T�R�"�a���j�U������53��68���2��6�6q�5.p�J75�2��J6�7�ǒ��(nU��A�5$ɼ�ɝ9|�J76��5�l�����63��77ֽ�578��60�a�54��J��4,I�81I�50'���a�6$�87q�NVuD5�7l�J67I�,�R84a( 7� �(6m�6�(7L���(Z�(9��64q�7��D0�F�8RTS���5�'SVM�BS�CTO��M��DLP鶊 %�NN�A�NNM4��EkXTQF[�88�IAB��J6 ��-׺3�6OPIQS�END��H�7PC�T�641(7%�C�PRe���@��ETmS�GGZ�FSG���0�X9�GSVH�M�SVS��.P�FG�TUq�GDѶSL�Ma�6H�G2��CP��W׍��_�_�_ 
oo.o@oRodovo�o �o�o�o�o�o�o *<N`r��� ������&�8� J�\�n���������ȏ ڏ����"�4�F�X� j�|�������ğ֟� ����0�B�T�f�x� ��������ү���� �,�>�P�b�t����� ����ο����(� :�L�^�pςϔϦϸ� ������ ��$�6�H� Z�l�~ߐߢߴ����� ����� �2�D�V�h� z������������ 
��.�@�R�d�v��� ������������ *<N`r��� ����&8 J\n����� ���/"/4/F/X/�j/|/�/  H59AD�!�!�5N�#R78	4�%5�*8N0�D�#ATU�4�$�54�4�&E4�#VC9AT�#CLI�4<4�RI5;UIF�*6�;CM�5|6:ST!Y�D�%HUl56UT<4�NR�Tl55�*R5�2%:�@�+S0U<4D�SB�:PL�T�#L;IC�:DOC�DLD�CSUf;9�:OR�SRf;8�*R86t�T�%0�:EIO�:�R54�*r@%:ES1E�T5$;J7$;�@��*MAS�T�#PRkXY�<7�*OCE:@P�:0�*P�,3UZ[J6�,53�JH�\�LCH5ZO3LJ5�0�:MHG�JPS4KM3LMC�;`[=5�;MDSWfkd[;OPd[MPRE:@�UZMAEN�,�\0.�*PCMe;0�kPX�:`�[51;5�l�50:PRS�JR�5tKJ69UZFR�DU:FREQ�*MuC�jS�LH93�*�SNBAf;�[SL]CU:SHL%KM�\@%:SPP�\2�\�2�:HTC�:TMqI�:� �JTPA�JoTPTXv�EL�k�50�K8�+� �*J�95�:TUTe[9�5UZUEV�JUE�C5ZUFRU:VC��VCO�JVIP�:CSC��CSGt�:c@I�)WEB�:7HTT�:R6�<�l0��CGԛIG��oIPGS�RC�:�DGd[H79:H.�LR76�;8Tk��n:R85u�66��7�KR#|�@��d�������0�53{6U8|2u\6%|6�;]5�;J75��25|T[J6��7t[�0u� T����5}u{5�MĬ:�]9�;J76�L䬱5�r@�;63�[7�7�+575�8u[60��54�Ӽ�pU�Y4%��K81�K5�˴0��6�L87�:N�VDe{7�J67�LkR84����Ҡ*U�6[6d�7��R����t�9�,64�;7�īD0��F��RTuS�{5d�SVME;;BSUJCTO�:b@��JDLPUJ���KNMNu{NN5���4�*�EXT5�FCm88.%:IAB��J��<tkc}6D�OPI5��SEND6ZH��P[CT��64��7�J�CPR�{�R UZE�TSGZ
SG�K��e̔�9��SVH�JSVSJ� 
�GTU�{GD5JS+LM�K6ԋGbpv�CP�:W�[�(�� �����
//./ @/R/d/v/�/�/�/�/ �/�/�/??*?<?N? `?r?�?�?�?�?�?�? �?OO&O8OJO\OnO �O�O�O�O�O�O�O�O _"_4_F_X_j_|_�_ �_�_�_�_�_�_oo 0oBoTofoxo�o�o�o �o�o�o�o,> Pbt����� ����(�:�L�^� p���������ʏ܏�  ��$�6�H�Z�l�~� ������Ɵ؟����  �2�D�V�h�z����� ��¯ԯ���
��.� @�R�d�v��������� п�����*�<�N� `�rτϖϨϺ����� ����&�8�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|�� ������������� 0�B�T�f�x������� ��������,> Pbt����� ��(:L^ p�������  //$/6/H/Z/l/~/��-� STD~�$LANG�$ �)�/�/�/??'?9? K?]?o?�?�?�?�?�? �?�?�?O#O5OGOYO kO}O�O�O�O�O�O�O �O__1_C_U_g_y_ �_�_�_�_�_�_�_	o o-o?oQocouo�o�o �o�o�o�o�o) ;M_q���� �����%�7�I��[�RBTq�� OPTN��������ҏ �����,�>�P�b� t���������Ο��� ��(�:�L�^�p��� ������ʯܯ� ���$�6�H�Z�l�~���DPN�$����̿޿� ��&�8�J�\�nπ� �Ϥ϶���������� "�4�F�X�j�|ߎߠ� ���ڑ(���� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v������� *<N`r� ������// &/8/J/\/n/�/�/�/ �/�/�/�/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $ 6HZl~��� ����� �2�D� V�h�z�������ԏ ���
��.�@�R�d� v���������П�������6�H�Z�l��~���99���$�FEAT_ADD ?	������ɠ  	 ��ү�����,�>� P�b�t���������ο ����(�:�L�^� pςϔϦϸ�������  ��$�6�H�Z�l�~� �ߢߴ����������  �2�D�V�h�z��� ����������
��.� @�R�d�v��������� ������*<N `r������ �&8J\n �������� /"/4/F/X/j/|/�/ �/�/�/�/�/�/?? 0?B?T?f?x?�?�?�? �?�?�?�?OO,O>O PObOtO�O�O�O�O�O �O�O__(_:_L_^_ p_�_�_�_�_�_�_�_  oo$o6oHoZolo~o�o�o�o��DEMO� r��   ���m�o0' 9f]o���� ����,�#�5�b� Y�k���������ŏ� ���(��1�^�U�g� �������������� $��-�Z�Q�c����� ��������� �� )�V�M�_��������� ���ݿ���%�R� I�[ψ�ϑϫϵ��� ������!�N�E�W� ��{ߍߧ߱������� ���J�A�S��w� ������������ �F�=�O�|�s����� ��������B 9Kxo���� ���>5G tk}����� /�/:/1/C/p/g/ y/�/�/�/�/�/ ?�/ 	?6?-???l?c?u?�? �?�?�?�?�?�?O2O )O;OhO_OqO�O�O�O �O�O�O�O_._%_7_ d_[_m_�_�_�_�_�_ �_�_�_*o!o3o`oWo io�o�o�o�o�o�o�o �o&/\Se �������"� �+�X�O�a�{����� �����ߏ���'� T�K�]�w��������� �۟���#�P�G� Y�s�}��������ׯ ����L�C�U�o� y�������ܿӿ�� 	��H�?�Q�k�uϢ� �ϫ���������� D�;�M�g�qߞߕߧ� ������
���@�7� I�c�m�������� ������<�3�E�_� i������������� ��8/A[e� ������� 4+=Wa��� �����/0/'/ 9/S/]/�/�/�/�/�/ �/�/�/�/,?#?5?O? Y?�?}?�?�?�?�?�? �?�?(OO1OKOUO�O yO�O�O�O�O�O�O�O $__-_G_Q_~_u_�_ �_�_�_�_�_�_ oo )oCoMozoqo�o�o�o �o�o�o�o%? Ivm���� ����!�;�E�r� i�{�������ޏՏ� ���7�A�n�e�w� ������ڟџ��� �3�=�j�a�s����� ��֯ͯ߯���/� 9�f�]�o�������ҿ ɿۿ����+�5�b� Y�kϘϏϡ������� ����'�1�^�U�g� �ߋߝ������� ��� 	�#�-�Z�Q�c��� ������������� )�V�M�_��������� ��������%R I[����� ���!NEW �{������ �//J/A/S/�/w/ �/�/�/�/�/�/�/? ?F?=?O?|?s?�?�? �?�?�?�?�?OOBO 9OKOxOoO�O�O�O�O �O�O�O__>_5_G_ t_k_}_�_�_�_�_�_ �_oo:o1oCopogo yo�o�o�o�o�o�o�o 	6-?lcu� �������2� )�;�h�_�q������� ԏˏݏ���.�%�7� d�[�m�������Пǟ ٟ���*�!�3�`�W� i�������̯ïկ� ��&��/�\�S�e��� ����ȿ��ѿ���"� �+�X�O�aώυϗ� �ϻ���������'� T�K�]ߊ߁ߓ��߷� ��������#�P�G�Y��}������  ������ +�=�O�a�s������� ��������'9 K]o����� ���#5GY k}������ �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-???Q?c?u?�?�? �?�?�?�?�?OO)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_I_ [_m__�_�_�_�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o /ASew� �������� +�=�O�a�s������� ��͏ߏ���'�9� K�]�o���������ɟ ۟����#�5�G�Y� k�}�������ůׯ� ����1�C�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ���������)� ;�M�_�q߃ߕߧ߹� ��������%�7�I� [�m��������� �����!�3�E�W�i� {��������������� /ASew� ������ +=Oas��� ����//'/9/ K/]/o/�/�/�/�/�/ �/�/�/?#?5?G?Y? k?}?�?�?�?�?�?�? �?OO1OCOUOgOyO �O�O�O�O�O�O�O	_ _-_?_Q_c_u_�_�_ �_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o|�o�i  �h �a�o/ASe w������� ��+�=�O�a�s��� ������͏ߏ��� '�9�K�]�o������� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� �)�;�M�_�q߃ߕ� �߹���������%� 7�I�[�m����� ���������!�3�E� W�i�{����������� ����/ASe w������� +=Oas� ������// '/9/K/]/o/�/�/�/ �/�/�/�/�/?#?5? G?Y?k?}?�?�?�?�? �?�?�?OO1OCOUO gOyO�O�O�O�O�O�O �O	__-_?_Q_c_u_ �_�_�_�_�_�_�_o o)o;oMo_oqo�o�o �o�o�o�o�o% 7I[m��� �����!�3�E� W�i�{�������ÏՏ �����/�A�S�e� w���������џ��� ��+�=�O�a�s��� ������ͯ߯��� '�9�K�]�o������� ��ɿۿ����#�5� G�Y�k�}Ϗϡϳ��� ��������1�C�U� g�yߋߝ߯������� ��	��-�?�Q�c�u� ������������ �)�;�M�_�q����� ����������% 7I[m��� ����!3E Wi{����� ��////A/S/e/ w/�/�/�/�/�/�/�/ ??+?=?O?a?s?�? �?�?�?�?�?�?OO 'O9OKO]OoO�O�O�O �O�O�O�O�O_#_5_ G_Y_k_}_�_�_�_�_ �_�_�_oo1oCoUo goyo�o�o�o�o�o�a�`�h�o!3 EWi{���� �����/�A�S� e�w���������я� ����+�=�O�a�s� ��������͟ߟ�� �'�9�K�]�o����� ����ɯۯ����#� 5�G�Y�k�}������� ſ׿�����1�C� U�g�yϋϝϯ����� ����	��-�?�Q�c� u߇ߙ߽߫������� ��)�;�M�_�q�� ������������ %�7�I�[�m������ ����������!3 EWi{���� ���/AS ew������ �//+/=/O/a/s/ �/�/�/�/�/�/�/? ?'?9?K?]?o?�?�? �?�?�?�?�?�?O#O 5OGOYOkO}O�O�O�O �O�O�O�O__1_C_ U_g_y_�_�_�_�_�_ �_�_	oo-o?oQoco uo�o�o�o�o�o�o�o );M_q� �������� %�7�I�[�m������ ��Ǐُ����!�3� E�W�i�{�������ß ՟�����/�A�S� e�w���������ѯ� ����+�=�O�a�s� ��������Ϳ߿�� �'�9�K�]�oρϓ� �Ϸ����������#� 5�G�Y�k�}ߏߡ߳� ����������1�C� U�g�y������������$FEAT_�DEMOIN  ����������INDEX
������ILECO�MP s���K����A��SETUP2 �tK�U�� � N ��>�_AP2BCK 1uK�?  �)���"��%������N��� ���>��b��o �'�K��� �:L�p��� 5�Y�}�$/� H/�l/~//�/1/�/ �/g/�/�/ ?2?�/V? �/z?	?�?�???�?c? �?
O�?.O�?ROdO�? �OO�O�OMO�OqO_ �O_<_�O`_�O�_�_ %_�_I_�_�__o�_ 8oJo�_no�_�o!o�o �oWo�o{o"�oF �oj|�/�� e����+�T�� x������=�ҏa��� ���,���P�b�񏆟����9�����Z���P�� 2��
SY�SSPOT.SV�矓�*�TEMy*4�]� %]����n����?�ԯ�� r����EAL ����˯`�k����� �,�>�P���	�g�=��LSCH��¿Կi�l� ����"�4πF�X�����ߘ���IAO������p�k�!� ��*�<�N�`��� ��~g�*.VR ��>R� %* ��{�0�����3�PC@�����FR6:�����1��%�0�TX��Y���F�x������k��*.F>�J���%!	������	��-��STM��b�����N��	���H O�s��(:��GIF�juV������JPG Y�u�/�0/B/F5�JSH�q/��#�St//
Java?Script�/�CSS��/u�!?�-Cascad�ing Styl�e Sheets�!?s�AZ*.B�IN �/��FR�5:\d5�?#)A�utoZone �.bin fil9eM?\9DATk?}?��7�1 O�?�2dat��?��ARGNAM�E.DO��x \@lO*O�!�D�OYO�@�DISP�0�O�� �D�O�O�A#Q1_�O��VGN�/	_�߰_k��]%BU: s�ervo gun��_g_y_o�_2o��LD�_co��PRE�SS�_o$o�ol��%�Rg press J@a�oso�o�o�o>	�Pb�on���#P�/�*�j�C{%�ddistd@u���@��Xtx����TROK��"�4�ɏl��fbckupk�~���%����I�L��)TW?LOGVAR�*��<�џl�`%�Qtwloe�v�����,���P��Xq��� �AG���>�ӯn�o� ��z�����2���V���Xq����hBT_KL00=ᮿy,�����q� �vatun �util忮�TP�EINS.XML�ψO:\(�2_�AC�ustom To�olbari��PASSWORD(_~
^FRS:\���k�PPasswo�rd ConfiYg���	S"PA'_�FߕB��0��� %�TbZ`f�agnosiRO'ݬ�I�[ڻ�z�x��!��bWPAT�0���:�8�P���PS�pot App OProc���������T���������#���G���X�}� ���0�����f����� 1��U��yr �>�b�	�- �Qc���� L�p/��;/� _/�p/�/$/�/H/�/ �/~/?�/7?I?�/m?��/�? ?�?�?��$�FILE_DGB�CK 1u����0��� < ��UMM?ARY.DG�?\OMD:ODO���D� Summ�aryEO�[CONS"�:OO/A�O�OWA}�sole ���O��TPACCNľO#_%_H_SET�P Accoun�tin�O
�S�6:�IPKDMP.ZIP|_��
�_�_TE�dPExcepti�o\o�\0@MEMCHECK>_�O3OTo��AMemory� D��i(i�=)?aRIPE�O-o�?o�occ%�a �Packet L��O�e���b�aS�T>��o�o�o�o %�bSt��|	FTP�o�C��_g�Amment� TBD��gx���)ETHERNE&�a$�d�WAEthern�`��ura�_��qDCSVRF�����ms�� ver?ify alϋe��\���DIFF�ޏď֏k��c �di�ffm�!�a��CHG01b�I�[��oqX���#�!���2柀͟ߟt���'���3pj�Q�c��� ��|���VTRN��G.LS$�կ�|�zga<� Ope��r�a \A�tic���q|)VDEV@�i�W�i���ms�Vis��Devgice����IM��AG�_ڿ쿁��d��Imag$ϱ�UMPɰESȿ]�\������Y@Up��es� List	�*��p�FLEXEVEANZ�a�sό�oqO� UIF Ev�q��o�c|��)T?D:GUN1L�e�xw��ceGun�� file~�e����2�����ߐ��1�C���3[�m��������T�EQU?IP1.TX��������equip�3����N)
P�SRBWLD.C	M��x�������@�PS_ROBOWSEL�xLP�I��z�����|�Net�/IP�a�ߵ����)� GRAPHICS4D�����%4D� Graphic�s F�����x�bGIG�o��>bfGigE�Ȳ�n���bSM��/�*/ag�/E�mail�4�&�,bSHADOW�&///�/)�Sha�dow Chan�gO�f ��bRCMERR�/�/�/�6?ec� CFG _Error�tO ��/ �*�sC?MSGLIB.?? '?�?�5xr)�H�?�u0)�)�0ZD��O�?:OagZD��ad�?i<%�)�,@IRDG_REPORW�O1OCO�%iR��s �Repor+� ��;�bPRCS�W�@�O�O�OH_�BS�pot App �process 9l��`��LJ�V଀t_)_;_EMe%�`_���^�Rs!NOT�I���_�_Lo��N?otific��iO>���x)�|o�o��ēo�oC��� �o�oB��o(�oL�o p��5�Yk  ��$�6��Z��~� �w���C�؏g���� ��2���V������� ��Q��u�
���� @�ϟd�󟈯��)��� M��q������<�N� ݯr����%���̿[� ���&ϵ�J�ٿn� ��Ϥ�3�����i��� ��"߱��X���|�� �߲�A���e��߉ߛ� 0��T�f��ߊ��� =����s����,�>� ��b�����'���K� ��������:��3 p���#��Y� }��H�l~ �1�U���  /�D/V/�z/	/�/�-/?/�/�(�$FI�LE_FRSPRT  ��� ����(�MDONLY 1�u5�  
 ���R_VDAEX?TP.ZZZ�/�/�h?Ul6%NO� Back fi�le B?�e| n/�?X?�?�/�?#Oh/ GO�?kO}OO�O0O�O �OfO�O�O_1_�OU_ �Oy__�_�_>_�_b_ �_	o�_-o�_Qoco�_ �oo�o�oLo�opo �o;�o_�o�� $�H��~���7�I��$VISBC�K 8
1/3*.V�DJ����FR:�\c�ION\DA�TA\��r��Vision VD�2�����0�>� (�b��s���'���K� ��򟁟���:�ɟ۟ p�������a�ʯY�� }���$���H�ׯl�~� ���1�ƿU�g�����  �2��V��z�	ϋ� ��?���c���
ߙ�.����R����ψ��*LU�I_CONFIG7 v5v��۟ $ q�%6{ 5����� �2�D�R���|xz�|���� ����j���	��-�?� ��P�u���������T� ����);��_ q����P�� %7�[m ���L���/ !/3/�W/i/{/�/�/ �/H/�/�/�/??/? �/S?e?w?�?�?2?�? �?�?�?OO�?=OOO aOsO�O�O.O�O�O�O �O__�O9_K_]_o_ �_�_*_�_�_�_�_�_ o�_5oGoYoko}o�o &o�o�o�o�o�o�o 1CUgy�"� ������-�?� Q�c�u��������Ϗ �󏊏�)�;�M�_� q��������˟ݟ� ���%�7�I�[�m�� ������ǯٯ믂�� !�3�E�W�i� ����� ��ÿտ�~���/� A�S��dωϛϭϿ� ��h�����+�=�O� ��s߅ߗߩ߻���d� ����'�9�K���o� �������`����� �#�5�G���k�}���������V�xR�obot Spe?ed 20%�� �$6HV�  �xO\�$FL�UI_DATA �w�����V�~RESULT 3x���  �T��/wizard�/guided/�steps/Expertk�� "4FXj|�����Conti�nue with{ G� ance� ��//1/C/U/g/�y/�/�/�/ ]-�^��)0 ��_��/�/���ps�/9?K?]?o?�?�? �?�?�?�?�?�?�_� &O8OJO\OnO�O�O�O �O�O�O�O�O^�/�/tB_<6rip�  "?�_�_�_�_�_�_�_ oo*o<oNoOro�o �o�o�o�o�o�o &8J\_-_w��1?� Time?US/DSTd� ��"�4�F�X�j�|�������Enabl�ԏ���
��.��@�R�d�v�������]�/������v24�<�N�`�r��� ������̯ޯ𯯏�� &�8�J�\�n������� ��ȿڿ�����ϟ��C�	7��RegionϐϢϴ����π����� �2�D߳America|_ ~ߐߢߴ���������@� �2�D�/V�y��,ώ��b��ditorU�������,��>�P�b�t������ �Touch Pa�nel �� (recommen� )������!3E@Wi{��^�n����������accesm�7I[m�������Zl�Connect �to Network�1/C/U/g/y/ �/�/�/�/�/�/�/b腘���:? �!���Introduct|Ϗ?�?�?�? �?�?�?OO1OCO^o gOyO�O�O�O�O�O�O��O	__-_?_Q_  n$?n_�_
�aO�_�_ �_�_oo0oBoTofo xo�o�o[O�o�o�o�o ,>Pbt�D��qP�_xZ�_ ��_�!�3�E�W�i� {�������ÏՏ珦o ��/�A�S�e�w��� ������џ����� �:��a�s������� ��ͯ߯���'�9� ��J�o���������ɿ ۿ����#�5�G�� h�*���N��������� ����1�C�U�g�y� �ߝ߮���������	� �-�?�Q�c�u��� XϺ�|������)� ;�M�_�q��������� ��������%7I [m����� �����0���i {������� ////A/ e/w/�/ �/�/�/�/�/�/?? +?=?�^? �?�?X/ �?�?�?�?OO'O9O KO]OoO�O�OR/�O�O �O�O�O_#_5_G_Y_ k_}_�_N?�?r?�_�_ �?oo1oCoUogoyo �o�o�o�o�o�o�O	 -?Qcu�� �����_�_�_� 8��__�q��������� ˏݏ���%�7��o [�m��������ǟٟ ����!�3���� (���L���ïկ��� ��/�A�S�e�w��� H�����ѿ����� +�=�O�a�sυϗ�V� h�z��Ϟ���'�9� K�]�o߁ߓߥ߷��� �ߚ����#�5�G�Y� k�}���������� �Ϻ���.���U�g�y� ��������������	 -��>cu�� �����) ;��\��B��� ���//%/7/I/ [/m//�/��/�/�/ �/�/?!?3?E?W?i? {?�?L�?p�?��? OO/OAOSOeOwO�O �O�O�O�O�O�/__ +_=_O_a_s_�_�_�_ �_�_�_�? o�?$o�? �_]ooo�o�o�o�o�o �o�o�o#5�OY k}������ ���1��_R�ov� ��L����ӏ���	� �-�?�Q�c�u���F ����ϟ����)� ;�M�_�q���B���f� ��گ����%�7�I� [�m��������ǿٿ �����!�3�E�W�i� {ύϟϱ����ϔ�ޯ ���,��S�e�w߉� �߭߿��������� +��O�a�s���� ����������'��� ��
��~�@ߥ����� ������#5GY k}<����� �1CUgy �J�\�n�����	/ /-/?/Q/c/u/�/�/ �/�/�/��/??)? ;?M?_?q?�?�?�?�? �?�?���"O�IO [OmOO�O�O�O�O�O �O�O_!_�/2_W_i_ {_�_�_�_�_�_�_�_ oo/o�?PoOto6O �o�o�o�o�o�o +=Oas��o� ������'�9� K�]�o���@o��doƏ �o����#�5�G�Y� k�}�������şן� ����1�C�U�g�y� ��������ӯ������ �ڏܯQ�c�u����� ����Ͽ����)� �M�_�qσϕϧϹ� ��������%��F� �j�|�@ϣߵ����� �����!�3�E�W�i� {�:ϟ���������� ��/�A�S�e�w�6� ��Zߤ������� +=Oas��� �����'9 K]o����� ������� /��G/Y/ k/}/�/�/�/�/�/�/ �/??�C?U?g?y? �?�?�?�?�?�?�?	O O���/rO4/�O �O�O�O�O�O__)_ ;_M___q_0?�_�_�_ �_�_�_oo%o7oIo [omoo>OPObO�o�O �o�o!3EWi {�����_�� ��/�A�S�e�w��� ������я�o�o�o� �o=�O�a�s������� ��͟ߟ����&� K�]�o���������ɯ ۯ����#��D�� h�*�������ſ׿� ����1�C�U�g�y� ���ϯ���������	� �-�?�Q�c�u�4��� X���|�������)� ;�M�_�q����� �������%�7�I� [�m������������ ��������EWi {������� ��ASew� ������// ��:/��^/p/4�/�/ �/�/�/�/??'?9? K?]?o?.�?�?�?�? �?�?�?O#O5OGOYO kO*/t/N/�O�O�/�O �O__1_C_U_g_y_ �_�_�_�_�?�_�_	o o-o?oQocouo�o�o �o�o|O�O�O�o�O ;M_q���� ������_7�I� [�m��������Ǐُ �����o�o�of� (������ß՟��� ��/�A�S�e�$��� ������ѯ����� +�=�O�a�s�2�D�V� ��z�߿���'�9� K�]�oρϓϥϷ�v� �������#�5�G�Y� k�}ߏߡ߳��߄��� ��
�̿1�C�U�g�y� ������������	� ���?�Q�c�u����� ������������ 8��\���� ���%7I [m~����� ��/!/3/E/W/i/ (�/L�/p�/�/�/ ??/?A?S?e?w?�? �?�?�?~�?�?OO +O=OOOaOsO�O�O�O �Oz/�O�/ _�/�O9_ K_]_o_�_�_�_�_�_ �_�_�_o�?5oGoYo ko}o�o�o�o�o�o�o �o�O.�ORd(o �������	� �-�?�Q�c�"o���� ����Ϗ����)� ;�M�_�hB���� xݟ���%�7�I� [�m��������t�ٯ ����!�3�E�W�i� {�������p�����޿ �ʟ/�A�S�e�wω� �ϭϿ��������Ư +�=�O�a�s߅ߗߩ� ���������¿Կ� ��Z�ρ������ �������#�5�G�Y� �}������������� ��1CUg&� 8�J�n����	 -?Qcu�� �j����//)/ ;/M/_/q/�/�/�/�/ x���/�%?7?I? [?m??�?�?�?�?�? �?�?�O3OEOWOiO {O�O�O�O�O�O�O�O _�/,_�/P_?w_�_ �_�_�_�_�_�_oo +o=oOoaor_�o�o�o �o�o�o�o'9 K]_~@_�d_� ����#�5�G�Y� k�}�������ro׏� ����1�C�U�g�y� ������nП���� ��-�?�Q�c�u����� ����ϯ���ď)� ;�M�_�q��������� ˿ݿ����"��F� X��ϑϣϵ����� �����!�3�E�W�� {ߍߟ߱��������� ��/�A�S��\�6� ���l��������� +�=�O�a�s������� h�������'9 K]o���d�� ������#5GY k}������ ���/1/C/U/g/y/ �/�/�/�/�/�/�/� ���N?u?�?�? �?�?�?�?�?OO)O ;OMO/qO�O�O�O�O �O�O�O__%_7_I_ [_?,?>?�_b?�_�_ �_�_o!o3oEoWoio {o�o�o^O�o�o�o�o /ASew� ��l_~_�_��_� +�=�O�a�s������� ��͏ߏ�o�'�9� K�]�o���������ɟ ۟���� ��D�� k�}�������ůׯ� ����1�C�U�f�y� ��������ӿ���	� �-�?�Q��r�4��� X�����������)� ;�M�_�q߃ߕߧ�f� ��������%�7�I� [�m����b���� ��Ϭ�!�3�E�W�i� {��������������� ��/ASew� �������� ��:Ls��� ����//'/9/ K/
o/�/�/�/�/�/ �/�/�/?#?5?G? P*t?�?`�?�?�? �?OO1OCOUOgOyO �O�O\/�O�O�O�O	_ _-_?_Q_c_u_�_�_ X?�?|?�_�_�?o)o ;oMo_oqo�o�o�o�o �o�o�o�O%7I [m����� ��_�_�_�_B�oi� {�������ÏՏ��� ��/�A� e�w��� ������џ����� +�=�O�� �2���V� ��ͯ߯���'�9� K�]�o�����R���ɿ ۿ����#�5�G�Y� k�}Ϗϡ�`�r����� ����1�C�U�g�y� �ߝ߯������ߤ��� �-�?�Q�c�u��� ������������� 8���_�q��������� ������%7I Z�m����� ��!3E�f (��L������ ////A/S/e/w/�/ �/Z�/�/�/�/?? +?=?O?a?s?�?�?V �?z�?��?O'O9O KO]OoO�O�O�O�O�O �O�O�/_#_5_G_Y_ k_}_�_�_�_�_�_�_ �?
o�?.o@o_goyo �o�o�o�o�o�o�o	 -?�Ocu�� �������)� ;��_Dooh���To�� ˏݏ���%�7�I� [�m����P��ǟٟ ����!�3�E�W�i� {���L���p���䯦� ��/�A�S�e�w��� ������ѿ㿢��� +�=�O�a�sυϗϩ� �����Ϟ���¯ԯ6� ��]�o߁ߓߥ߷��� �������#�5���Y� k�}���������� ����1�C���&� ��J߯���������	 -?Qcu�F� �����) ;M_q��T�f� x����//%/7/I/ [/m//�/�/�/�/�/ ��/?!?3?E?W?i? {?�?�?�?�?�?�?� O�,O�SOeOwO�O �O�O�O�O�O�O__ +_=_NOa_s_�_�_�_ �_�_�_�_oo'o9o �?ZoO~o@O�o�o�o �o�o�o#5GY k}�N_���� ���1�C�U�g�y� ��Jo��noЏ�o��	� �-�?�Q�c�u����� ����ϟ០��)� ;�M�_�q��������� ˯ݯ������"�4��� [�m��������ǿٿ ����!�3��W�i� {ύϟϱ��������� ��/��8��\߆� H��߿��������� +�=�O�a�s��Dϩ� ����������'�9� K�]�o���@ߊ�d߮� ������#5GY k}������� �1CUgy ����������� ��*/��Q/c/u/�/�/ �/�/�/�/�/??)? �M?_?q?�?�?�?�? �?�?�?OO%O7O� //|O>/�O�O�O�O �O�O_!_3_E_W_i_ {_:?�_�_�_�_�_�_ oo/oAoSoeowo�o HOZOlO�o�O�o +=Oas��� ���_���'�9� K�]�o���������ɏ ۏ�o���o ��oG�Y� k�}�������şן� ����1�B�U�g�y� ��������ӯ���	� �-��N��r�4��� ����Ͽ����)� ;�M�_�qσ�B��Ϲ� ��������%�7�I� [�m��>���b��߆� �����!�3�E�W�i� {����������� ��/�A�S�e�w��� �������������� (��Oas��� ����'�� K]o����� ���/#/��, P/z/<�/�/�/�/�/ �/??1?C?U?g?y? 8�?�?�?�?�?�?	O O-O?OQOcOuO4/~/ X/�O�O�/�O__)_ ;_M___q_�_�_�_�_ �_�?�_oo%o7oIo [omoo�o�o�o�o�O �O�O�O�OEWi {������� ���_A�S�e�w��� ������я����� +��o�op�2���� ��͟ߟ���'�9� K�]�o�.�������ɯ ۯ����#�5�G�Y� k�}�<�N�`�¿��� ����1�C�U�g�y� �ϝϯ��π�����	� �-�?�Q�c�u߇ߙ� �߽��ߎ��߲��ֿ ;�M�_�q����� ��������%�6�I� [�m������������ ����!��B�f (������� /ASew6� ������// +/=/O/a/s/2�/V �/z|/�/??'?9? K?]?o?�?�?�?�?�? ��?�?O#O5OGOYO kO}O�O�O�O�O�/�O �/
__�?C_U_g_y_ �_�_�_�_�_�_�_	o o�??oQocouo�o�o �o�o�o�o�o�O  _�ODn0_��� �����%�7�I� [�m�,o������Ǐُ ����!�3�E�W�i� (rL�������� ��/�A�S�e�w��� ������~������ +�=�O�a�s������� ��z��������ԟ9� K�]�oρϓϥϷ��� �������Я5�G�Y� k�}ߏߡ߳������� ����޿��d�&� ������������	� �-�?�Q�c�"߇��� ����������) ;M_q0�B�T� x���%7I [m���t�� ��/!/3/E/W/i/ {/�/�/�/�/��/� ?�/?A?S?e?w?�? �?�?�?�?�?�?OO *?=OOOaOsO�O�O�O �O�O�O�O__�/6_ �/Z_?�_�_�_�_�_ �_�_�_o#o5oGoYo ko*O�o�o�o�o�o�o �o1CUg&_ �J_�n_p��	� �-�?�Q�c�u����� ����|o����)� ;�M�_�q��������� xڟ����ԏ7�I� [�m��������ǯٯ ����Ώ3�E�W�i� {�������ÿտ��� �ʟ��8�b�$��� �ϭϿ��������� +�=�O�a� ��ߗߩ� ����������'�9� K�]��f�@ϊ��v� �������#�5�G�Y� k�}�������r����� ��1CUgy ���n���� ��-?Qcu�� �����/��)/ ;/M/_/q/�/�/�/�/ �/�/�/??��� X??�?�?�?�?�? �?�?O!O3OEOWO/ {O�O�O�O�O�O�O�O __/_A_S_e_$?6? H?�_l?�_�_�_oo +o=oOoaoso�o�o�o hO�o�o�o'9 K]o����v_ ��_��_#�5�G�Y� k�}�������ŏ׏� ����1�C�U�g�y� ��������ӟ���	� �*��N��u����� ����ϯ����)� ;�M�_���������� ˿ݿ���%�7�I� [��|�>���b�d��� �����!�3�E�W�i� {ߍߟ߱�p������� ��/�A�S�e�w�� ���l��������� +�=�O�a�s������� ����������'9 K]o����� ��������,V �}������ �//1/C/U/y/ �/�/�/�/�/�/�/	? ?-???Q?Z4~? �?j�?�?�?OO)O ;OMO_OqO�O�O�Of/ �O�O�O__%_7_I_ [_m__�_�_b?t?�? �?�_�?!o3oEoWoio {o�o�o�o�o�o�o�o �O/ASew� ��������_ �_�_L�os������� ��͏ߏ���'�9� K�
o���������ɟ ۟����#�5�G�Y���*�<������$F�MR2_GRP �1y���� �C4  �B�c�	 c�x����E�� ���\��P]��Q�*.a<�Nȗl^D�M�D(�?&�x`�\��:�?>���8��(�A� � ��»BH�C�K  ܶ`�\��x
���@UUU0��UU(��i��>���
?��?>���>�1>��ff>H�9(�;�D���o;�ı�H���l���� ��+��O�b�ܯz� � Z߱ߜ���������� ��¿P��u���� �����������;� &�K�q�\������������`���_CFG {z˫T "���+=O��NO �˪F270�477 �� ���R�P
���RM_CHK?TYP  ��c�pӠՠ����ROM� �_MIN� c����� ��X��SS�B{�� v�c���1��TP_DEF�_OW  c�|ӣFIRCOM� �W��UNC_SE�TUP  ˫������GENOVRD_DO��m�c-�THR�� d%d�_E�NBv �RA�VCģ|��  ��ߊ/���/�/r�q�/�/�� �y/ ?�/B?T?�/c?�/	1�Z!O�1�ˬ rc����<� �r��?�?�?�?(OfԖ@ް�1XO�5rO]ݬ&�oFBȉ�oB���9�O�?�7O8O_B�O_I_KG�^_�_�_c��&��O�O�_�RSMTģ�h)נ� MDLE�$HOSTCs2�˩� �m�k 	KhKkKo2c�{o`�e�o�o �o�o�o_��o/AS�e�o�p	ano?nymous������ Jo\ono K���o������ɏ ����#�5�X�� �}�������ş�� 0�B�D�1�x�U�g�y� �������ӯ���	� ,�b�t�Q�c�u����� �������L�)� ;�M�_Ϧ�pϕϧϹ� �����6��%�7�I� [ߢ���ƿؿ�ϴ�� �����!�3�z�W�i� {�������
����� ��/�v߈ߚ�H��� ���߿��������� +=Oa����� ����8�J�\�n� K�������� ��/#/5/X� �}/�/�/�/�/ 0BD/1?xU?g?y? �?�?��?�?�?�?? Ob/?OQOcOuO�O�_~-aENT 1�9i?�  P!O�O `  �O_�O (_�OL__p_3_|_W_ �_�_�_�_�_o�_6o �_Zoo/o�oSo�owo �o�o�o�o�o2�oV z=�a��� ����@��L�'� u���]�����⏥�� ɏ*����`�#���G����k�QUICC�0����!172o.19.��11ܟ@ė�����S�ƕ2U��1�C���!ROU�TER�����25�4̯t�PCJO�G��Я�9��68�.0.10ΟÓC�AMPRTE�!�!�5�1>�l�S�RT�p���� !S�oftware �Operator? Panel��2��3ϩDNAME �!�J!UB10200RBT0���HS_CFG 2���I ��Auto-st�arted�$FTP�/��?O�� D?�-�?�Q�c߰?�� �߽߫�����t��� )�;�M��.�Ϸ��Ϧ� ���Ͻ��� ��$��� H�Z�l�~�����5���@������ �'r��Strt Vis Prt���q�� ���������� %7I[~ ~� ����38J\ �p]/��/�/�/�/ �/t/�/�/?#?F/G? �/k?}?�?�?�?�]? 	�8((�8/:?'O n/KO]OoO�O�OZ?�O �O�O�OO�O�O5_G_ Y_k_}_`�)_�?�?�_ _/O�_o0oBoTo_ xo�o�o�o�o�_eo�o ,>P�_�_�_ �_�o�o���� (��oL�^�p������ 9�ʏ܏� ��$�k }�l��������Ɵ ؟꟱�� �2�D�V� y���u�����¯ԯ��<�_ERR ��T���PDUSI�Z  ��^�����>2�WRD �?�� !�  gues  ��r���������̿C��SCDMNGRPw 3����g� $}�׃��!����K %	�P01.m�8�� �  I  
��A�మ�	�?� �������(i���u�R�u��Y�  2 W n��@���E��"��>�g�������������8m������5 ����  ��A�����s����[��s���i�m�)�����YH�3�5 (5  �d=�O�a�s��h}䃦(�09� �=��������:�%�^���d�g���M� "��K������*��__GROU����_  ޲	���4�ڶ��A�QUPD'  ��A���TY  ��S�VG ��ֺn�< �?�S�B �������݃������ "4FXj|� ������ 0BTf}�����TTP_AUTH� 2����!i?Pendanط!.�y���C!!KAREL:*!/*/<-�KCQ/a/s/I �VISION SETK��/�/B'�/�/  ?�/G??0?}?T?���P�v?�?�?�4�CTRL �������
9ЮFFF�9E3�?b�FR�S:DEFAUL�T/LFANU�C Web Server�@+§� �Z�l��<�O�O�O�O��O�O �WR_CONFIG � �� o/O�IA_�CHKCMB 3�� �L�
 ���4�?�_�U [�c��R�R��P�Q�S�� d��_��t��_�_zVo �_�_�_�_�o�W�o�o �o/o�oSoeowo�o�o E[I�o�+ =O����\�� ������Ï��K� �o���������a�w� e���ğ#�5�G�Y�k� �+����x�ן��� ��ɯ߯ͯg�,��� ������ӯ}������ �?�Q�c�u���1�Gϼ5�YRDEBU��� g]P��E��������~L_DEL �g[��< �A���8F��UVELBa_s] l�����/�#�5�_� Y�;�ɿ_�������� B�0�*���N��r�� ������������� &�8�J�\�������W ��{������^L Fj/����  ���BT fx���s/��/ �//,/z/h/b/'? �/K?�/�/�/�/.?? ?�?:?�?^?p?�?�?��?�?�?�O}�FOBoJ 3����'@	P]L�3���O�OYOp�O5_G_^ <>� `߂_�Sn_�_�_�_�_ �_�_o*ooLo�O Ae�O%_�o�o�o�o�o e_;oAo9[ ]o�����Oo ao(��o�op�����W� i�ʏ܏'���� �K�1�S���g�y��� ��#�5�G�����D�V� �+�����i���џׯ ��߯���'�)�;� ]������п�}�� �*��N�`�rϽ��� ��k��ϳϵ������ ���Mߧ�����ݿ?� �����߯���"�4�� E�g�i�?�u���� ���������{ߍߟ� �����A������ ��S�)�/�7eK ]����=�O� (s���^p�E� ������/ //A/o/U/w/�/� �/5� ?2?D?? ?z?�?��/�/�/�/ �?�?�?O1OO)OKO MO�/�/�/Y?k?�O_ �?�O<_N__�?�O�_ YO�_�_�_�_�_�_�_�o;o�O�O�n�$I�A_GRP 3������a?� L*U*o8Lo�o�d	 @�o�o 
o�o@"4V� j|�����'� ��N�0�R�����x����̏������ 
� 0&X)Q'P� �  �C��  R��[�B�D��N��X���E����&TB�^N�Z���  B��������+ꮒ�d�4%�ʜZq��N��d�z��Si��&Tj��N�2��S�B�� _� ?�u�X�j��������8į���  p�$�p��K�l� |>� `���8���̿���� ����J�k�>�`ϒ�pxϚ�����[�
���E^�  к� g���� �d!�%�&�8�
� �=�)�$Ce�ntral Pl?ane Ck9�z� �ߞ߰���������
� �.�@�R�d�v��� ��zo�Ͼ�����o� P�q�D�f���z����� ��������
L. @b�v���� �3(Z0�� �������/� �<//`/C/U/�/y/ �/�/�/�/�/�/&?	? ?Y;�5Gi�?y� �?�?�?�?�?!OO%O WO=OOOqO�O�O�O�O �O�O�O�O"XD�߀�s_rL�^�p�o_  �e�e�_�_�_�_o o 2oDoVohozo�o�o�o��o�o�o�o��%S�$�IA_LCFG ���e�J%P�4�\Q/��ks�<6�<�s,gs�S��qur64�� }FsOG 3�R{'
 l�%S!!� 3�%�Q�c�
�i����� ��Ïj�Տ����/� ֏A�e�w�����B��� џ�������=�O� a�s��������ͯ߯ ����'�9�K��]� ��������^�ɿ�����;}NET ��R}_'_^�(�UM_�CHK  j�c�\s
��ELB<�ϥ�FOBJ�ϥ�x�q�Ϧ�PAIR�ϛ ��WTߥ�O�TF ��e�� �D/  BH  ?=���A Dtһ3�R{ �}puP�aQ P?�j�L?�����߯�� "�\�����y��� `�����6�H���-� ?���u�������^� ����������);�� �����j���v�GqSETUP ��R{`QTRA1K�Y 
 �	
��@ G�i�S�OG�k} �����/�/dO/n,� ?2�\P�/�/�*2�.gP��\ UQ  ��\ Fb � 
_�$b�PZ\ ���q\ 	�MQ� $\ �qbp�"��b 	8
�$�q�op]\P� ��C4?8?8op�,C46�a\P�b F0�\P�qNPB1�qe�8NP�0=b �.pٯ4� ��Q�b 0�6� :�4��4�!� "\ s�b NP?\ b ��8`pgPpb TH@@b0 q�,1F۰�� mb �0-
@�b #�$ZA0)�p�kQ� 6��e� &�0��Ȳb '`0YP*b (J\ �b �b nA|�DV�@e\P�b +� �� �b �p>��m�O�O_G �� \&C/e/?_%_G_ u_�_e_�_�_�_�_�_ o�_o;o!oCoqo�n  _~o�oVo�o�o �o �o6.P~\n ������o�
� D��L�z���j��� ��ʏ����
�@�&� 8�v�\�&�t������� ؟������4�V� ��b�t���̯��ԯ� ����J��R����� p���ȿ�������� �F�,�>�`�bϯϼ��@�� ��WTP:|Х��
 ����20M�F@ ߷�Z��d��XI�UU@ؕ�2^������� ;�M�_�q߃ߕߧ߹� f������'�%�7�I� ��m��������� ����!�3�E�W�i� {���:���������� �ASew� ���l�� +=Oa/��� �����//'/9/�K/],��B_CHK?CMB 3��Ʌ!Ŵ�'!�/m/�% &@�&~%�%�(PC?�"���?�?�?*5�? D?V?h?z??O�7@OVO DO�?�OOO&O8OJO �O
_�O�OW_�O�O�O �O�O�_�_�_F_oj_ |_�_�_�_\oro`o�_ �oo0oBoTofo& �os�o�o�o ���b'���� ��x���|��ۏ:� L�^�p���,�B�0�ʏ ��� ��$�6��������2DEBUG �=�^���J����n�����/�L ��;�$wϙ��ìELB?"=������� �!ҟ����x�� m�������߿ٿ�� ����!�3�E�Wϥϓ� ��R߱�v�������� Y�G�A��e�*�ߛ� �߿�����ߺ���� =�O�a�s�����n� �������'�u�c� ]�"��F�������� )�5�Yk }������� 1C�y>/�,�FOBJ 3��;���P,� ���/�//�/�/�/�. <��1?<3? ??m?S?u?�?�?�?�?�?�?7/�5r/�/]O oO�ODO�O�O�O?�? �O�?�O
___@_n_ T_v_�_�?O�_4O�O o1oCoooyo�o�O �_�_�_�_�o�o�o 0(JL�_�_�_ Xojo���o�;�M� ��o���X������ ��֏؏��:��� ��,���ǟٟ���� �!�l�B�H��@�b� d�v���Ư��ί��V� h�/����w�����^� p�ѿ�.������ $�R�8�Zψ�nπϢ� ��*�<�N���¿K�]� �2ߓߥ�p������ ��������.�0�B� d��������"߄�� �1���U�g�y��ߚ� ��r���������� &T������F� �����);�� LnpF|��� �������� �/�/H�/�/�/ �/Z0/6?/>?l?R? d?�?�?�?�?�?D/V/�/N�$IB_GR�P 3�����LA� L��%�?�?yO�D	 @ aO�O�O�?�O�O�O�O _7__+_M__a_�_ �_�_�_�_�_�_o3o To'oIo{o]o�o�o�oO 
 0�(�!� �   �c/C�  u�
p�g��e��b�s�a�SE�4v�$�h^�a>	u��  Bjpeu�IxPt�]r�p4h�oy| q��a�pMz7ti��v�$x���a�a�t�u�  �/�b�t$���Z�=��O���s�����  �rӏ�o�o��� |��E��M�{��� o���ß��˟������A�'�I�w���[��
��E^�  �б� r�n� d�"d � S012SSW�01���k���i�m$�Centra�l Plane Ck�)�;�M�_�q� ��������˿ݿ�� �%�7�I�[�)O[�m� �ϑ��O���� ���� G�)�[�}�c�qߓ��� �߹��������C�%� 7�Y��m������� ��	��j����[�>�� b�t����������� ��E(:{^� �����Ώ�� ���R(�B�f� ����/�� / N/0/R/�/j/|/�/�/2�(D�r�� Hïկ 2?����1w<LELE u?�?�?�?�?�?�?�? OO)O;OMO_OqO�O�O�O���#�$IB�_HAND 3��E� 
�p4�c�/_�(_^_ A_S_�_w_�_�_�_�_ f��_�!_�_Bo%o7o Io[o�oo�o�o�o�o �_o!o�oP3EW i������ ��^�A���e�w� �������я��+� ����O���s���Ɵ ����͟ߟ �'�9�� ���]�������ԯ�� ɯۯ�.�5�G��v� �k��������ſ� ���<�C�U�'τ�� yϺϝϯ�������� 	�?�J�c�5ߒ�)߇� �߽߫�����"��� M�_�q�C������ ��������0��%�[��m��BLCFG ]�[  t�K��  ܯ�S6l�!��,�����
��6J<����U4}��OG 3�\ l�#!�Oew P9��N���� �=Oas �������/ '/9/K/�]/�/�/�/ �/^/�/�/�/?#?�/ 5?Y?k?}?�?6?�?�? �?�?�?�?O1OCOUO~�MNET ���� <{� ?��aK�OaO�BPAIRw 3�[ � �T T P�J X�_1_C__ g_y_J\�OM___�_�_ �_�_o*o�_�_oro �o�oYoko�o�oAoSo �o&8J�� �oi����"��4��O��SETUP� ���T ��J�K�p
 �	
~�@�O�O��ȋ�� ���Џ�$�E��:�@l�N�������~�J��K��ڟ���2>؞  ��py�_  ��pFJ V�
_:�6 Z�p-G���p�6��$�p:��P��J 	RZ�
B�:��]K�t�ِ�������������U�a�K��q��K���( ����ި ���=J  ����U��J ]��J�:��ّ6�U"�psJ  ?�p�J V���)��pJ n�]�]�f��  ��@�?�imJ M�a��J �#N���i�)��ԲJ %6�Ѡ/J &��K���J '������*J (�p�J �dJ ű|���eK�e�J +*�=��J ������.�@�<R�`� �4��� ������|Ϟ����ϼ� ������J�k�:�\� ��xߚ�����w���� ���)�W�5�G��k� ������������� %�S���?�a���9��� ����������!O p?a�}��� }���/]; Moq����� �#/	/+/Y/�E/g/ �/?/�/�/�/�/�/? ??U?;?E?g?�?�? �?�?�?O�!�Β] sBWTP�@�~K
 �Ot�����u�YD��wOM�qΑd n�VBhȠH�q�q�H͗2�CKO]OoO_�O�O �O�O�O�O�O_�_5_ G_Y_k_}_�_�_No�_ �_�_�_oo1oCo�o goyo�o�o�o�o�o�o �	-?Qcu "�������� �ď;�M�_�q����� ����f�ݏ���%� 7�I���m���������*@C_3D_CF�G �j���G~"_�AZ�_CALIB 3�m���?�?��x��~#0��  ��D�V�9�z�]�o������Կ�ɿ
��  �&�O�B�\Ͻ?��ү �������������9� �]�o�Rߓ�v߈��� ������z��5�(�B� k�ϸϒ�������� ������C�U�8�y� \�n���������`��� (Q|��x� �������) ;_BT�x� �F�/�/7/b �^//�/��/�/�/ �/�/�/!??E?W?:? {?^?p?�?,/�?�?�? �?OH/j/DOeOwO�? �O�O�O�O�O�O_�O +_=_ _a_D_V_�_O �_�_�_�_�_.OPO*o Ko]ox_�o�ovo�o�o �o�o�o#G* <}�_����� o6o�1�C�^�y� \�������ӏ��ȏ	� �-�?�"�c������ ����������0�)� D�V�_�B�����x��� �����ү�%��I� ğm�h�r�������� ���*�<�E�(�i� {�^ϟςϔ��ϸ��� ���/ߪ�(�N�w�j� ��ƿؿ�������"� +�� �a�D���z� ���������'��� 4�]�P�j������ߺ� �������G* k}`����� ���C6Py ���������� �-//Q/c/F/�/j/ |/�/�/�/�/n ?)? ?6?_?���?�?�? �/�?�?�?O�?OIO ,OmOObO�O�O�O�O T?�O___E_p?�? l_�_�_�O�_�_�_�_ �_�_/ooSoeoHo�o lo~o�o:_�o�o�o V_x_Rs��o� �������9� K�.�o�R�d��� ���ďΏ����et�$I�C_AZ_CON�F �����:��epTdxJ� ep_�<ep�+�MEMBR ;3�:� H��������џ��� ����9�7�a�C��� �����ɯǯ�ӯ� �9��Y�W���c��� ��ɿ������1� /�Y�;�y�wϡσ��� ������	��1��Q� O�y�[ߙߗ��ߣ����*�PROG 3�:� ��ew0�B� o�f�x�������� �����5�,�>�k�b� t����������������1(�SCHE�D 3�:�  HRepG�J�dep
�����Voxel ?Sched1ev����2��.�!3v�4Se���5��/�6��N/�7+/=/�/B�8s/�/�/�9�/(�/&?���	0?? o?:>�T?f?x?�
 �?�?�?�R�?�?O ��,O>OPO��tO �O�O�*&�O�O�O� r&__(_��&L_^_ p_�6�_�_�_K? �_>o	o�?-o�oQo�? uo�o�o#O�o�okO ^)�OM�q�O ���C_�6���_�%�~�I��_m�Ə�^3 o���ُco��V�!��
`PACE 3�� �������� 	 ��D��  E	� D�e���B� �C���� ��,��  �?aG���:�� @���̟ޟ���ѯ 8�J�\�n��������� ȯگ��z��"�4�F� X�j�������]�Ŀֿ �����0�����f� xϊϜϮ�������� ���,�>�P�b�t߆� 0�&���������� X�:�L�	�p���� ������� ��$�6� H�Z�l�������L�� ������ �DV hz������ ��.@Rdv ���i/���/ /*/</�/�/r/�/�/ �/�/�/?�/?�?&? 8?J?\?n?�?�?<O���LST 3���4 6O�;NO4O�O�O�O�O �O_�O_V_5_G_�_ k_}_�_�_�_�_�_�_ �_oo1oCoUogo�o �o�o�o�o�o�o*	�`?Q�uZJD�P_CONF ѯ��>�D�
K�d h�0�>�rE�0Ez�0�;� ?8Q�@7��́{�`A=���uSCHED 3����
�D�eadlock Prevent�p 8�������� ͏��ڏ����9�,� F�o�b�|�����ɟğ Ο�����"�0�Y�L� f�������ů��ү�� ��1�$�>�g�Z�t� ����������q\�n� ȿ1�$�>�g�Z�tϊ� ���ϼ���������� (�Q�D�^߇�zߔ߽� �������� �)��6� _�R�l������ ������� �I�<�V� ��ω�p������� E8R{n �������
 A<Fwr|� ����/�/=/ 0/J/s/f/�/�/�/�/ �/�/�/?'?����? o?b?|?�?�?�?�?�? �?�?O"O0OYOLOfO �O�O�O�O�O�O�O�O _1_$_>_g_Z_t_�_ �_�_�_�_�_�_�_o (oQoDo^o�ozo�o�o 0?B?�o�o
$M @Z�v���� �����I�D�N� �z�������ُ̏� ���E�8�R�{�n� ���������ڟ��
� �A�<�e��o�oD��� ��ѯ̯֯���*� 8�a�T�n�������Ϳ ��ڿ����9�,�F� o�b�|ϒϘ������� �����"�0�Y�L�f� �߂ߜ��߸�����n� ������U�H�b��~� �������������  �Q�L�V��������� ��������
$M @Z�v���� ���IDN z��(���� /
//2/@/i/\/v/ �/�/�/�/�/�/?�/ ?A?4?N?w?j?�?�? �?�?�?�?OOO*O 8OaOTOnO�O�O�O�O �O�O_�O_9_�� �*_�_�_�_�_�_�_ �_�_o"o(oYoTo^o �o�o�o�o�o�o�o�o ,UHb�~ ��������  �Q�L�V��������� ���T_f_�ҏ�:� H�q�d�~�������ݟ П��� �I�<�V� �r�������ٯԯޯ �
��2�@�i�\�v� ������տȿ������A�4�N�w���$�IC_DP_SI�D 3�������� � u�jƻ����� ���0�'�9�f�]�o� �ߓ��߷��������� ,�#�5�b�Y�k��� �����������(�� 1�^�U�g��������� ��������$-Z Qc}����� �� )VM_ y������� //%/R/I/[/u// �/�/�/�/�/�/?? !?N?E?W?q?{?�?�? �?�?�?�?OOOJO AOSOmOwO�O�O�O�O �O�O___F_=_O_ i_s_�_�_�_�_�_�_ oooBo9oKoeooo �o�o�o�o�o�o�o >5Gak�� �������:� 1�C�]�g�������ʏ ��ӏ ���	�6�-�?� Y�c�������Ɵ��ϟ ����2�)�;�U�_� ������¯��˯��� �.�%�7�Q�[���� ������ǿ�����*� !�3�M�Wτ�{ύϺ� ����������&��/� I�S߀�w߉߶߭߿� ������"��+�E�O� |�s��������� ����'�A�K�x�o� �������������� #=Gtk}� ����� 9Cpgy��� ���/	//5/?/�l/c/u'�$IC_�DP_ZID 3߳����!� d / u/�/�/�/?
??I? @?R?l?v?�?�?�?�? �?�?OOOEO<ONO hOrO�O�O�O�O�O�O ___A_8_J_d_n_ �_�_�_�_�_�_o�_ o=o4oFo`ojo�o�o �o�o�o�o�o9 0B\f���� �����5�,�>� X�b�������ŏ��Ώ ����1�(�:�T�^� ����������ʟ���  �-�$�6�P�Z���~� ������Ư����)�  �2�L�V���z����� ��¿����%��.� H�R��vψϵϬϾ� ������!��*�D�N��{�rߑ*DL_CP�U_PCT�Є�B��  �� B�;MU��MIN�ܱ!� >jQ� GN�R_IOERR � �ӯ%�#ICD_BG ��)���-iicmedCbg��G���\�d���(�i3��W��h�iisv2���V���~�'��� �.�o ��s���L�^����:�~��)ud1:����*�DEF 1��%p�#�-��.����buf.txtp���_CF�q��s�� y��������
�3��d� p�����ZSTATE �3��%!�
 �p�"������/���>/-/@b/Q/�/u/�/���/ �/�/�/�/"??F?��5?v?e?�?�?�?�? �?�
�?OO7O&O[OJOO��mO�O�O�O �O�O�O_��	_J_ 9_n_]_�_�_�_�Z�_ �_�_o�_/ooSo��	Ao�oqo�o�o�o�o �o�oC2gV��
��!����NPT_S_IM_DO����'�tL_SCR�N�� ���T�PMODNTOL�H��_�_PRTY�'���x�VIS��E�NBH���_F_FRCVR���	<x���M  ̋z�	���RSMPRG�ɏ�����$IO�LNK 1�,� Y�������Ο�����|�MASTE������OSLAVE� �,�2�RAM�CACHE"�Z�O_AUTO�e�|��|�UOP��v�CMT_OP����0����YCLc���, _A_SG 1�|��p�)�;�M�_�q��� ������˿ݿ���\s���NUM��0��
x�IPa�s�RTRY_CNů��D�O_UPD�ӗ���1 x�����,�� ��Ϙ ��P_MEMBERS 3�|]s� $����v�� ٪��RCA_ACC �2��  S�X@��r6#�z�*�pqn���ߒ֗գ�P�BUF�001 2��=� R@u2  �u2R`u3��3�R��Ԡ���������S����S u4���4S@���S��!���S���Tw uF��FT Y�0�T��T@�TH�T��TX�U����U T����U��U �U�UU�U�V �V��MV0�V`�� �VH�SV����W��Wh��W0�W��X tr� @�X u?��?�X0�XI%�  W%�P��P �PH�UP�P�Q��Qh�UQ0�Q��Q@�QH�UQ�QX�R��R����2�������#�5� G�Y�k�}������ ��������1�C�U��g�y�����������3����    	    !��)�� 1��9��
$H��Q��"$`  ho q o B$�o R$�o "$�  �� �� $��� $�� "$�  �� �$�� �  $� � *$(/0 z$8/0
$HO0QO0B$`  ho0$xo0"4�  ��0z$ ��0
$��0Z$��0�j$� �$PԹ�2���{ <!�	J0W  <p#D&A)�P��HIS��±{ �܎� 2021�-08-11vC ��&@)�&@yDU yD(yD0yD8yDE@yDHyD��$BX�E �A&A�O�O�O_ _rS
�``H�BpO�OP�O�O�O#C`UThUTEpUTxUT��%A�UTU�UT�UT�UT�q�;  l2&@�UT�l�Q&@S	:Y09H_ Z_l_~_�_�_�_�_�_ �\&@l2�Pnj`b (o�S@oRodovo�o�o��o�o�je�Pb�PSj7 6o$6H Zlr�Pt���nj6�� ��$� 6�lZ�l��Px���jj5��ʏ܏� � �$�6�l�Z�l�#C;I ��JO\O������̟ޟ �O���"�4�F�4_F_ ����ůׯ����"� �_F�ooy������� ��ӿ���	��o�o�o�c�uχϙ� :� �	 3 >�� ! ,���� ���ϴ��W�E�W� iߟ�D��߱���D��� ����/�A�S��w� @����v���������s�9�K�]���� ��\��o�����3E�� C��@��@l�$��� @)�n1D�^2K�- ?QcQ�c���� �@%@-@ 5@=@E@M@ U@�@�@l2@ )�@1�:ϕ�� ���//%/7/I/ �q/�/�/�/�/�/ �/�/??%?��M? _?q?�?�?�?�?�?�? �?O��)O;OMO_O qO�O�O�O�O�O�O ��__)_;_M___q_��_�_�_�_w`�I_�CFG 2Õ� H
Cycl�e Timew�Busyw�Idl�b�dmi�nt
qUp|�f�aRead�gDow�h�o{��q�cCount>�a	Num �b�c��tz}wRq`�P�ROG�bĕ�� �)/sof�tpart/ge�nlink?cu�rrent=me�nupage,1133,�����'�|w`�SDT_�ISOLC  ��	� n�sR�_USED  a���bJ23_DSPo_ENB�� ��?INC ŏ�w�o�A��?= =�̟�<#�
n��:�o ���w��E�K�JOB�pC䩃�U���pGRO�UP 1�a�~��d< �{p��v��M�?Qv  �GUN:�{͟ Q�%�7�I�� m������w5�wd<��ǟ��۟� ��e�^�p���A������ʿܿ�� �|�IN_�AUTO����PO�SREg���KANJI_MASK�V���KARELMO�N Ǖ�wy �����������s�{�J�sȱw��w'�|Bϼ�KCL_L��NUM��\�$KE�YLOGGING��� ������pLA�NGUAGE �����DEFAULT ��6�LD�aɱyA��r>��q��G�aʬ�z
r�Vdm ���)�w'� _ � 
�w�wy6�D�;��
~�(UT1:\��� �������� ����0�=�O�a�x��c�ϴ�x��N_D?ISP �ʏx��� ����OCT�OL9�Dz�pj�A��!GBOOK ��d��q���[ :e��������� �r�	�	�A����Gd��?_BUFF 2��a� U2 u�ZE��w�� /�
/7/./@/m/d/ v/�/�/�/�/�/�/�/�?3?���pDCS �����A����e��?�?�?�?J4IO ;2��� �`O�`�p�
OO,O>ORO bOtO�O�O�O�O�O�O �O__*_:_L_^_r_��_�_�_�_�5ER_ITM^�d��o%o 7oIo[omoo�o�o�o �o�o�o�o!3E�Wi{�RSEVte����VTYP^��o����}>�R�STz�H5SCRN�_FL 2��=�{?{�������Ï�Տ��TP���^��rNGNAMpU�3�����UPS��SGI0�G���V��_LOADPRO�G %�z%C�C�0����MA�INT_�?��  (%��ퟘ� ۟���8�#�\�G��� k�������گů��� "��F�X�C�|�g��� ��Ŀ���ӿ��	� B�-�f�Qϊ�uϮ��� ���������,��P� ;�t߆�qߪߕ��߹� �����(��L�7�p����XUALRMN3UMb��u�0���\�a�d� 5 � p��C����K������_G�RP 2�K �ؚ	�q�  ��E��>�j� U�g���y8�������� ����)M8q� f������ %I[>j� ������!/3/ /W/B/{/^/p/�/�/ �/�/�/?�//??S? 6?H?�?t?�?�?�?�? �?O�?+OO OaOLO �OpO�O�O�O�O�O_ �O�O9_$_]_H_�_�_�v_�_�_�_��DBG?DEF ���������_�P_LDXD�ISAA��{Y���E�MO_AP;�E {?�{
 a X�dovo�o�o�o�o�o��o��FRQ_CF�G ���cAM X�@�)sX�<��d%�lQ�op�����9��*�p/�r **: �rX��xCX��� ���E�<�N�{��_ �夏`��ˏ���،,(y�"�X��M�4� q�X�������˟��� ��%��I�[�B�� ������u�k���� �2�)�;�M�_����� ��������ѿ��,� g�P�7�Iφ�mϪϑ� ���������(�:�!��^�E߂ߔߊ�ISCg 1�Si�p �� ��9�o���_"��F� X�?�|��ߋ�_����������_MSTR� �Sk
`�SC/D 1�Sm���`� ���o����������� ��&J5nY ~������ �41jU�y �����/�0/ /T/?/x/c/�/�/�/ �/�/�/�/??>?)? N?t?_?�?�?�?�?�? �?O�?O:O%O^OIO �OmO�O�O�O�O�O _��O$__H_3_l_�M�Kq� �}_�LoTARM
r�w�R �p�_��T�Rxq_DO �ܙ_.�p�������U9oy��3ohoWo�o{o�_$M�METPU(`y��(�qNDSP?_ADCOL�e#a�mCMNT�o/��b�FNp�gFST�LI,w� ݀ �~�S!b� c�eP�OSCFMw~PgRPM
�yST�`{1�>� 4@y�<#�
���+� 9��9�;�M���q��� ŏ������ݏ�1���%�g�I�[������aS�ING_CHK � /$MODA�Q�R߱ۧ[�Y~әDEV 	>��	MC:�ڒHOSIZE(` ��וTASK %>��%$123456�789 x���՗T�RIG 2�>� l>�%}�د��Ư ����=��2�s��FZ�YPE���֓�EM_INF 1���W��`)�AT&FV0E0�x��)ױE0V�1&A3&B1&�D2&S0&C1�S0=޽)ATZ�C�*�HG�o���c���&�A���ς������!� տF���� �/Ϡ�S��������� �����B�T�;�x�+� =߮�a�s߅����� ,�c�P����A��� �������������� ��^������k� �� �6���� l1C��y� !/��D/�h/O/ �/�/Q�/u��� ?�@?R?�/v?)/�?�U?�?�?�?�?�^ON�ITORhpG ?��   	EOXEC1cS7B2=H3=H4=H5=H��?FU7=H8=H9cS8B �"�D<B�DHB�DTB�D `B�DlB�DxB�D�B�DP�B�D�B�C2�H2�HU2�H2�H2�H2�HU2�H2�H2	X2X�3�H3�H3HBבR�bSV 1�Ļ� (����?����g �:�ϻ�5˿Ǫؾ篚�z���G�1YOOb�_D�2H��%cION_DBG� ���  +��`l�`m�tjdk }�~wg�k`��k`�t�0N  � -��`�wk���p��-ud1�1��o�o�o?qPL_NAME !��(p�!176�908 iB/7�00 E-SG �Ax�TRR2�Q 1���x�y�(q�p\ d�r u������� ��)�;�M�_�q����������ˏݏ��2 q�,�>�P�b�t�����������	���� 
��.�@�R�d�v��� ������Я����� *�<�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶��� �������"�4�F�X� j�|ߎߠ߲����������P<՟"�4�F�X� j�|����������$y��"�
�F��TP5�r��������� ������&8J \n�O�a���� ��"4FXj |������� //0/B/T/f/x/�/ �/�/�/�/�/�/?>� D�� C�� 22�Y  �G?Y=�RdC3+0x?�= n?�?�7,0=�]? O�?$O'4�PG@O6O HOZOxO~O�O�O�P;`h�O�L�RE	`*O�$_6_H_Q:�o�ALrh_z_�_�� 1B�`�Y?7��c�a�1s`�BM���B0$�RW�  �Z90��de
O +oOOoaoLo�opo�o }p�o�o%7 I[m���� ����!�3�E��� i�{�������ÏՏ� ���ԟA�S�e�w� ��������џ���� �+�=�O�a�s����� ����ͯ߯���'� 9�K�]�o��������� ɿۿ����#�5�G� Y�k�}Ϗϡϳ����� ������1�C�U�� yߋߝ߯��������� 	��-�?�_�U�}� 4������������� �1�C�U�g�y����� ����������	- ?Qcu���� ���)��M _q������ �//%/7/I/[/m/ �?�oX?�/�?�/�?�/ ?�?�/�oW?B?{?2O �O�O�?�?�?�?�?�? �OAO�O
_wO�O�OR_�d_�O�O�O�TA�  Yk?0_g<iZ_o &_�_~_�_�_�_�_�_�o� �$MRR_GRP 1�\@�3a;`*@nBj�5 ^B~Ha @D�  \a?�bcHa?� da�!�@2��Ez  ��a(�o  ;�	�ltb	 ��`L �`��qPrP�`X0w&��`� ��b�� K�e�K����b���K�jK���\f��_��/)�q?���Dv�f�Pq|a5C��Iۿ��5��6�����F{�q}�4�  �e`�f�ô�p��sb`k�����q��$	�`�R��rua��L_j_v�  �j@�KH��  ?�  �T��_�r�u	'� �� ��I� ��  �Uv:��È��È=��9�̅r@܏� �~Na�5Nb�"��wN�@^�  '�t�p@up?�p?
�@�p@�p��L��C�pB�pA�  EC�pB�p��7*@߼�D/�c�� �I���X`�l ����@�BP��M�4�qD�ea�^�I����m�����O� ��� ��[`���ѐ�  �r:��ef�*@0�?��ff'?�$��� !]@Y�k�q8p��^��>�R`pa�z=	  �����PAǳ�q�c�d�&�>Lր ѐ�hq;�~�;D�A g;�-�<���o�?? B&�7tb�Nc��P?fff�?�?&n�4D@�{����A
��� 7ؒi�udyde��bg ��RǨdC���<�'� `�K߄�oߨߺߥ���x��F�@����� >��_���1��-�� ������������4�� X�C�|�g�����=�������oU�y�H���ᙕF�,�A  3�` ?�����B����`i{��:�A��p)H:���w�B�a���	B-�AA�fY��C8���%� 3/����}�؂����2/�uč�Sâ�̩���D�^`;��
�P�����rD\Y�C��s3C��B�33BZPɱ�}� ���� A�333�̀���/��9�3�ٙ���_��Bm��A�33�/���0;� nffBd�p ���[
<pL����L��K3�ÜIĮIK��G�d��E1��3,L�4L��ʖIb� I-ߞ�G��_?���4LA�L�?��I���Ir�H#��?�?�8�\!�?�?OOqA{
?,O: KOTO�OxO�s�O�O�d�|�O�O J	)��O�OJ	��5_�OY_ D_: a/k_�_�_�_�_ �_�_�_"ooFo1ojo Uogo�o�o�o�n�!�o �o�o�E�@�od�'�_t� ?�� ���!��Bc����L�Z�O� L���3�>�KI�[�f�����Ï��ӏ����G뵐�ێD_�;$��o�Z���~�0����۟ƟCf���֟7��"(�!3f��;�����l�$��G��\�n��3�����3|������L�|3z	����D���E�w3����L�@:�p�^������P�	Pƾ�����B��� %��I�4�m�Xϑ�|ϰ0*������1� E �ϊ����7�"�[�� ����|߲ߠ������ߜ��
�<+J�� :~ ��4���|�j������� k 2� ��7C�����B�ne�C�Z n�@u:�L�@^�p�lڂ_����� �������$�p0T������8���
 � ������� #5GYk����oH稤���:��� @D���?��� � `?<�!��A�X����j�;�	l�ñ0s �,ñ d(,��G�N/���@|/�,��9�/�)�/@�/R�?�//?�$u��P?^8!7����  Р?�8!?�?	�9�?�? == O&K�)����BOLF9F&�jOxG�㿠O��'�O�L�A��c�O�O_ݦ��a/�9_�B)�~_ >��U�AECױ_�_�_�_�_o�_ �#c �!-o;g  �Q!:o�1[OHda���\qo�oo v��o�k�8�P�o�j>=#���9o+S_	�>L>"gb�!(�y@�o(�����P�?fff?>�?& �p�_����q���� $��D��v$�x�c� ���������Ϗ��8�>��� F�-� z�)������9���� ����:�%�^�I�[� �������ܯǯ �� �?3���Z���{�ٟ�� �ƿؿ�����#π��V�A�z�eϞω�����ip���ϖ��� �ʏu���F�1�j�U� gߠߋ��߯������ ��0�B�-�f�Q��u� �����������,� �P�;�t�_������� ��������:% 7p[���� � �6!ZE ~i������ � //D///h/z/e/ �/�/�/�/�/�/
?�/ ?@?+?d?O?�?s?�? �?�?�?�?O�?*OO NO9OrO]OoO�O�O�O �O�O�O_�O8_J_5_�n_Y_�_}W(������_�[�_�_�_
o �_.oo>o@oRo�ovo��o�o�o�o�o�l�P�rP&~E�"ԅ_V �X[�p���� ��� ��K�6�o� Z���~���^ ��D� ����=�+�a�O��� s�������ߟ͟��'�5�  2��[�m� �������ǯٯ�����J�/�A�S�e�w�ࢌխ�����
  ��������0�B� T�f�xϊϜϮ������"rۿ���}���$MR_CABL�E 2�x ���T<p@w@  /� ?�0��.�*��  ´�  BK�CGК�O4>�B���r�9bJ��`��Fr?g.D�Rۚ�+�~=��4  ��L��7pB���N�Yк^Ф�by ��_�n� ?D���(�bߑ�TH�L���\�Ъҋ�0^З�b�
��an�#}D�.�����@�-B!�x߾>�8� J�\�n���������� ��?����:�4�F�X� j����������ᚱ�q ^�^з�^Я6�^УJ��R�b�^��r��*��������� ������`��� �����@������ ����`�$� �)� /@�ĕ ʙ Ϡ���@*�  ����)���� ���M jDV� z������� I//f/@/R/�/v/�/ �/�/�/�/�/�/E??�b?<?N?�?r?�;CH  ��*�?OO+O�� �?XOjO|O���?����OM �����i�  ���ą%% 2�34567890	1�O�E �O_�A��U𚰠�������
 W�Nnot sent�
��1P�WuTES�TFECSALGR  eg��3�-Q�d�T2T
�T3��<p�����_�_�_���9UD1:\�maintena�nces.xml�oNo  >t����DEFAUL��ԑV�GRP 2��J  �����<���  �%1�st mecha�nical ch'eck ]�����a#��c�o4��1�W�$6HZl���cc�ontrolleAr�d��o�5�����"�4��qMX�m\���"8r�#b�x�w����̏ޏ��?�C�"�q�F�v��t����������q�C�a�poling fan��3��xc�8�J�\�n���ڃrC�`ge�b. battery��'  3����7�ȡϯ�e	'���� �2��D��q��grea�seH���f���-�p�����e���ҿ�����W�Supp�lyb�t������Q����ϖϨϺ��σq���cabl,ϥr���
�<�p�ߪe
 s�H�Z�l�~ߐߓ��q����~7����0�B�T�qOve�rhauU�{l���� x�p���e������������p$ ��@��8�?o��2���� ���������S��� w�L^p����� ��=$6H Z�~���� ��/ /oD/�� z/��/�/�/�/�/5/ 
?Y/k/@?�/d?v?�? �?�?�/�??1?OU? *O<ONO`OrO�?�O�? �?�OO�O__&_8_ �O\_�O�O�O�_�_�_ �_�_�_M_"oq_�_�_ jo|o�o�o�ooio�o 7o�o[o0BTfx �o���o�!�� �,�>��b����� ���Ώ����S�(� w���^����������� ʟ��=�O�$�s�H� Z�l�~���ߟ���� �9�� �2�D�V��� z�ɯۯ����Կ��� 
��k�@Ϗ�����i� �ϬϾ�����1��U� g�y�N�`�r߄ߖ��� M���߻�?��&�8� J�\�߀���߶���������"�����	� X2�_�q�����B ��������� ����J\,� ��t���� �FXj(:�� ����//���(, ���?� ; @�� ���/ �/�/��w/�/�/ ?���* ?** F�@ 0!.&� R/X?�j?|?>?�?�?�?�?�����:?�?*O<O NOOrO�O�O�O�? O fO�O__ZO�OJ_\_ n_�O�O�Oz_�_�_�_ �_o"o4oFo�_�_o �o�o�o�o�o�o�o�Ro3����J��!�Vt��  �~�56@+������ ��nC�F/���� N�`�������0���� ޏx�9��p����� ��˟����>��֟�� 6�H���l���X���� ٯ��N�����p�E�W� �{�ʯ��b��¿p� 6�Ϫ��Aϐ�e�(� ڿ��6�����pϪ�� V�+��Ϡ�N����ϗ� 6�p�����ߴ��� �߈�]���6���߷� z������N�#����� ���.�@�����|�� ������\�����T f����v�"� �l,�Pu< x���2��T )/;//_/��/F/� �/T//�/�/�/%?t/ I??�/l??�/�?T? �?�?:?O�?�?2O�? �?{OOTO�O O�O�O �O�O�OlOA_�O_w_ �O�_^_�_�_l_2_o �_�_z_�_o$oro�o `o�_�olo�o@o�o �o8Jo�o�Zl ��P��r4� Y� �\����d��ď r�8����C���g� *�܏��8���ӟr��� 	�X�-�🢟P���ğ ��8�r�ϯ�󯶯h� �į��_���8���� ��|�ʿܿ��P�%�Ŀ ��[Ϫ��BϐϢ�P� ��ϊ���^�p���� V�h�D��ϱ�Pߊ�$� �߼�n��.�S��w� >�P��߿��4����� V��=��@����H�����V���s�	 X`��/s�B �� ^�������v� � ��HZl *<��r��� /�� /V/h/&/8/��/�/�/�/�/�/��� �~�?�  @s� <7?I?[?�s�#?�?�?�?s��*�?** F�@ �!�&w0�/OO(O��?LO^OpO�O�� �����?�O�O�O�O�O _0_B_T_�O�O_�_ �_�__�_�_oo`_ r_�_&oto�o�oZo�o �o�o�o8oJo�o:L ^p2����o����s��$MR_HIST 2��%}�� 
 \&��$ 2345678901"�*���2!�9�����J�|� �ۏ�����ȏ5�G� Y��"�p�����j�ן �����ğ1��U�g� ���B�����x�寜� 	��ү?���c�u�,����s��pSKCFM�AP  �%��x2�qs������ONREL � s��ʱ�p��E�XCFENB��
8ȳ���FNC���JOGOVLIM���d�e���KEY���h��v�_PA�N����³�RUN�X�h���SFSPDTYP<�Ų��SIGN���T1�MOTZ����_�CE_GRP 2��%ʳ���y? f�s�Sߐ���z߻�r� ���ߨ����%�K�� o�&�h��\������� ���#�5��Y��c� ��v���j����������A��*SYS�TEM*�V9.�3*�6 D2/1�2/2021, ���p1��MTC�OM_CFG_T�    $�CNC_NO۰�$NORES_T�IME�OPW�ORKp ,� $2 BUSY>�p$SOP����T�
U�INT�P��NING�P�AUSED�MA��OPT_OUT�۰�_DISA�BLEIMA�GE   �_PREV_IyM� /INV_ �/RW�RDVAL.�SERP.wPS_�L_O��� $|�MLT�_RBT{�p$�PMC_EDT_�� NOALM��DUMMY1�94�[SL�CT� � �$OVSL� �$SDIHDE�X1��2�OF[F_"VR'N!D#" #''"(�G#CS_CT�V!$'^\_ZER��_SETUP��0r#NUMn$E�RRID  �
�&_S�*�!�!���ARMLOAD����$�$� � �'�"v0�&_yP�#�!MRR26�>� 0�!���RA� � d$CA?LIB_MO�!� /GEAR/82J8 � $SPR�� ��43<$R>0S�W0�4#ABC�_FLAG�D_�J2SEC� �23�6
�21SP����! P�4�=3��=CUR_�� R�5J#E3�V"�� f1 	$CScKP��9ELI�&9EJN�15AQ:LkE�QEkEaGEXT_A�Z�C�AELEV�DhVOCMPT�OL2DAXISI�NERTI�F�%1)@�%X�@�HP ��JZ�DSMGRS�T� 2DJGFL_�SC��@ �AS/PH_I�"<U � ;0RT� ��!�$S[PA_LE��!:PGRATIO��#4B{TDI�A)R2[3U<BDF��Q�LW�XVEL=AI�NR� RT_BL�� 	�Uf2*Q�T�W�W�UMECH�_��E#RTSA�_1��!� ER%A�2/eI��Q,-b3`_N�<eWb�U,cWa�"	ai�V��DH5PV`�
 0� $_I'!$L7SP!$P:PW8R�0:P!D15H �$BE��ENG@\P_AC�CE�Q� w!pIGRC_|P��T�A�#�zXP{�Bu�JO� $wQ@L1%vPATHyzwszw�3�PROCESS_���c�p�qbR:P�C^pp_M��9QD1D�q|R8RFW� � `
s�usr�xDE��� BNQwRO?PEE�r:P8��aAA�DEFLXq'af�_<0�PINY RBx�Y*��`ҮY{ �GAR@�� � ��M�OU�qNG�pO8�PlqńINC� bA :P��t/�@�f1��7ENClPLE�3�A�Ps�yINPOȉ�.�M�#+PNT|�S�UNT23_�R�8R\�LO�P8Rr�E aQ�|��P	dA4 N0�O�M��pA�MO.�� ��T�q���3CPERCH  �
c�"�ۗ�A�STO��֗��G�B���p$�p(CA�;�Lx�(C0�ɒ'GD�UP���z���TRK_U� PCAY�#5�f���YHs�������FA��@M�OM߂􂹡AMP�1�T�07ţ|s@���`�2�sS_BCKLSH_;��<������ ���1P�e���cECL�A��8�� ��CHK�������RTY_ST��a�Q0�`�U��_��#��_UM��C����q2Q�C�LMTF�0_L�`�C�U3)�E �A�3��6u<ŀ6x�0P���F����P�C��HORTM9O�v�CMC��@\p�wCN_K2N�L��#SF�a�V���a$�[Q���%պ�CAT�SH�#K2�t �۱%�%��%��)�@f�pPA��_P� ԣ;1Q��ϐ=A����ĵJG�0Tp�Uq�P�OG��gRTORQAUt��5��ʩ�O� 0�rgR�8�_W�����A�aW��cV��cV�I*^�Il�I�cFn I�B��!A�pVCp0e��T��1���p��RA���J� ���
�'@Df~SM�S'@MC�0sDLP!U�GRV]�`V��cV��c7�H_�#85�}p��COS���@��LN�����P  ��P����������2�1Z��Ŗ7�MY��0��TH��Q	THE{T0��NK23�c�{7S��CB�CB7SC@0AS�!���0��c��SB�c�N�GTS�C�C�1@��G���G������^�,02�U;�UQ��_�C�QNE��iqKѴ�I�X] oA�s��������LP!H��zT�zS��� �����z��#*�] V�V��`�V��V�V +V+V*+V*+V8)H����"�Z��(�H +H�+H+H*+H8)OJ�O�Oi9�O�UO�O +O+O+O*+OFz��9���D�SPBAL�ANCE_@,CLmE� H_sSP4a���TB��TB��PFULCXHBgGB��Aj{1�UTO_���ĵT1T2�I r2N��3�L��D�����@P_Pr�c��Tk�O�P|qG�INSEG3����REVV��0�D3IF��fi1KW�R1	��OBAQ��`���2"�L���?�LC�HWAR*�0�AB���c��@ ��e
�X��Pe��V��b�@
 
�R5��a&�7ROBϐCRC�e���  �VaEC�T�  H �$T�PðATU�SM���CdP_wIDXTfBTM`g�Ja�`gp0�MY4�i�6cDT�a DnF`EPT-�DEccxjq�UaFILEj���UaEXE[`��a�b�b�d7�@` @\Fa"pUPD&qo�>tPP_PXNd��e�q�d��i �PG�_C��@`, $SUBIa�U��_Ia�ٰMPWA�IG�Pҁ_wr��F�����D��RCVF�AIL_�p�dqR ��7pƃ���`�uĐz��L[sDBTBñBWD�vRES�UᰧuIGPAU�S_PR�A��TN1L���t�RT��QpOΐ%�ҁ|�T�2¹�HADOWð�S�p�*���R���3qDEFґ@` LF`�Pr�8ё3���UNI@�iā�qR�`7RN�_L���PSa D��PH_PKT7s�  �pTR1I��� �OU�r3a�̀�FIՂ �� $Ѐ�� 3}݀DBGLV�s?LOGSIZ��6�$Ѐ�qU4�:�D���3_T��QMM�@���7SEMI�RZ�CO|���VCHECK�p�Ł�PIN9q' 0��$�`t�8qQpT@KETĂC�+BU&Q��P�r?a� h �-� �~q�`����S;`OR~[sFORMAT�@�tCORD-�`�Ҵ9���UXW)���ޒLI�r?a $݀��SWI�P�Ãp�W7Ы��Z�LL�B?a� $3BA&�L�ON�a�p�A[�sPks���BA#J5q�&QϢ6զ�_KNOWœ�\ �U�a� D��Ѐ�DUS���'��V�4�Y3�Z3�LSq�PǑ�PL�ΰ ! n�ɡ" |���&���F��CRPOPj�~bm�}�Ij�RO �j��Ѷ`��BASE2?QJ7R��_Jt�!���@���b�t���� ���p�pAL_� h���A�BQB�{��D2�E���J3'�;� T~�PDCK_R���pǑCO���T°%B�K�]��>�C�_�q�  �\�@,�D_13�2]�D�������
Ӱ`_RTIA49�59��6�MOMENT@E�e�R�e�_Ӊ�Bxp�ADEӉ�RӉ�_�PU� NRjԶ�RӶ��_��a�'�?a � ��Q�0r��G�R�b� e$PIq��n�^�p�� ���\�������&`�W���V9�HIG w�9�yur���r�yu�p �p�����q��qyuSAMC@�A�sB��� C�yuĠ�1q�?PE ��Wq�����
�"!R)`>Ԉ�7�V	��IN��7�&��������yr����:GA�MM(Fa�\�GET��FIœ]��Æ�=
�@LIBR�a�yI�ړ$HI�`C_V��c`=B�E��b�A�� �LW� ���	����V��t�C�u�PER��Ro ��I_%��������6�����eӃ�փ;� ��@n� 1�I/M_SR�PDwS�Rq�t�PLE��٢���R(���M�MS�WFL�t��SCR�x10K@�``��3 !be&��?PEЙ�y)��ވ%PI3A�METHt1�� �u�"�P��R�`X<�� �ESRI�$B�3nR����_0��0;DC��$#2��209L�C�E5OOP���![1��N�!APP!%�F�� D@_5�4k5���@1:O�@��8�1�b3���@1-1�ԓ@�:u@��2RA��MG%����}P@`PQURK'AGR
`�b`�SA���@"a=E�cNO��C!�b��=@� ��>�P�\�J�K���X���H
�DOq�A� 9Q��{*����Ǒ��Ǒ`�;W7U�Cs� W�}M� � �YL,����d�U!b��WS1�Q貱c�_r�C$��aM_Wl@B�RK2�0�SG6M�p �[���W.цtT$���S%rmPM.A�b !���P� qWM`�$�0L�q`�M`�� Kb��Kb��Kb_��p� AN��n�[�7�X��	O��6�Z�emP�p�W ��2M�L� O�O�O�O�OVа1!�ƀ2�PL��_�  |~�x=@eٗvR� �v_�=@>��w�vX�}�(�szB!ǀa�{t�P��PMON_�QUG� " 8���QCOU�]�Q�THg@HO�RB�H�YS�ESʢB�U�E-�3B��O�# � ݀P+`�!RU�N_TO�S@O����$ P)���Cx�QZ @INDE�$ROGRA�P,��P}2K0NE_NOքƋ�IT��ـo�IN;FO�% j�������R�AOI�&{ (�0SLEQ��P*���*�_o�S]��' 4��EN�AByb��PTIOyN�	�ERVE��p����%�^�GCF/�( @6�J`6���+�� R�������STR\�_EDI�Tc�) �Z`�`K������E� NU���AUTYA�COPY��2���e@�M�N<�@�UPR�UT� C�N��O;UC��$G����vjQAPذCRE�*�r�PM�E�IZ��_RS�ET ۬��a��FRO����DЀ�䃅DSP_C`��$��TCH3@��TEM�PI�Ru@HST^��O_SN,�a!=W ALM_m"`�`���1q�d��ISs�d A/�B��襯������4�PRGAD�J��+ h~�X_�L0I��`ݶ�`ݶW۸P۸ ݶ��Ͱ�b�NEXT_CYCZˣȲNSc�,{P扱GOb��NYQ�EQ��W���n�צ!LA#e�۱`�����幠� �# IFlH�ʃNAK�%���_G#STATUx~p#��MAILI��w�� =�LAST���v@�ELԠ0�-� �ĩ~0EASI t�JRv�Z�%���n!W�2�� I���eQ0E��#��AB���@�Eπ��VѤ�BA!SRA�֙qU���R@$����RMP�R��� ���c���b��� wpB��c�.�p	c� 2-  �d��I��� H��*`q@�Q��t�u&DOU���z2@��P10�/1�GRIyD݁��BARSh֐}�u�m���O�pA0+ |�_��!	�����O�`r�1 �s ܀�pPOR����%�SRV��)l8�0�DI[@T_��PR�d���n�3l�4l�U5l�6l�7l�8P�қ�Fj/�2z�$VALU��0EI�����Fc�3� !p�fá���-H0AN/C�����0r�w?TOTAL_�ĊЖTPW[�I��iR�EGENg
|�sX��ؠ�E	�(�TR����g_S8��| �3V۱�������E���0G�v��(�0V_H��DA(s� .GS_YaA�bצS@`{AR(p22 ��gIG_�,SUP0��_��	C_��$cCMu0ne�DEp@i]�Ia@Z��n����ENHANC.�4�p
Ʃ���� *C�O��`F��a�MASK�#��OVR�$�0Dp���a��OVC����$�
0���5l���h֥���P�SLG�0�6 \ 9B��T�*dQ ��qS�RԧU\� ���%��$x���"?�>/�7 (�~��J�&YB��IL_MĎ�?0V��� �pTQ���& ���C�v�RVl;Cz=P_>0R@�3mM�9V1�:V1�;U2�;2�;3�;3�;4�;4�:����R���04F�QRINEIV�IB8`t4a@QhD2�dHZfF3dH3pH4dH4pH/��4zr8�����4F��@G=EQE=EPL��TOR,����D�US� �p.�8=d�PMC_FK�Z�	5�8Q7Q�G �M�p���TR�� �װ]r��PKE��H/NADDMQ!�T���YC�a0�T��NRTаSO!��TF�LQ�`��S��SREM�R@�T�����TahU���e�THPWD  ;�SSBM!	�?COLLAB�$ (� E���IO��a�:�NO]qFCAL�DDON�wp6Sn�d9 ,��FLH�>��$SYNFP�l�M�pC��� UP�_DLY�q:z�DGELA�`����Y��AD(q��QSK;IP+�; �(����OR��=Az�pP_ ����8w��H��Ow�� ]y��]y��\z��\z���\z��\z��\z��\z9���RA�< X�\+'MB�PNFGLIC���f�Ue�<���'NO_Hp�R�D�0SWI5��"R�A_PAЀG��=S ��ǨU��W���o�_�NGRLT �`������� � �t���T_J�qC���P��WEIGH��Jg4CHf���OR����6"OO= �vї�J  ��A�� ����OBr�r��J2T%��a>l�X��Th�_�IT/_�ʰ�R_��:!�Q$�RDC\)�b? ��R���XR��Z��SK�R�GEA�x�S��F�LG_Ы���� ER�[Q�BSPCn�3�U�M__�%32TH2�V��Q� 1> �S�ED��� @ D Ʃ����W2_P�m�S�!���L10_C��sFDB�! Aհ � h�`ҕ�y�U1����%��XAl�s�S � "z��	0C��C�N�B PT�DE�SIG��h�VL1br�1��1�10`཰71u1ƱPOS;11"qC lװ�Q0�"�Pi�scAT�PN��20UB���IND 0 %!��{�
U�����B�HOMEϲ�w�2�D��������Ϳ߿W 	w�3�Eπ�&�8�J�\Ϥax�4�Fϑϣϵ�������w�5�G��� ߠ2�D�V�pw�6�H�yߋߝ߯����� w�7�I����P,�>�P���8�Js��������� h�w�SS`"qK  ��x�� ���b��L TT���J&��IO"1��I.�vO�`_OP����D�󑎒�WEGAM# o�`}�@�D� N�e $DSB� GNA�C�`�C/����S232N��O ������P�0ICEt�,PE�r`#X�IT0/O�PB{`"FLOW�TR��#b0#�CU� ѠɁUXT�!#�ERFAC4k�PU� t0C ;CH"qP t�PIP�_q �Ɓ$FR?EEFROMH�#�Aِ�`�OQUPD�fP���PTf�E�X@p4!O FA0iP���C MF��PCK Q L�p{���� Mz-+�-E��$:!_d0�Q_DUMMY�q��qv�dCTRL/_ R'pf��4b�MA��FF0��S��PX����'GP��SECGF�p��`0P+!MOVE r8#s h_3Q �P�QR�O%�T$���c@�o@�bD� oS �`PO �+5�"�bV�qT7D �DS�c�X����r�DR
pU]12,�V�&EF�� ���s h"�'D'`;S$fALM�Pcbܑ @3INFJ7_H�AP{���@CB RYǃJ�!-!��%�$pcw�67RITR�>]RZ_OFFߢ�PAPA���»2�.n-�MNTwCMc�S��y�pjН3�#U� �693�5lP <0PF�84IECCad��HK�����!�l����COUz��G��ALA�2� �AU2��SPG&5	!2ZFD� R_ab-�Vw�!���3����M�Op ���7�STE���L(�RE�GDI_5!�Fd7�A# ��LTU��CVVrF�HP�B09��3�4�"A`EC�g�V 8\�MONq�@D�Vj`s ��R��U �RDI�B1� WR�UB1MSG�rEV�H�*�+�ED�`j��SSHAR�X <\���`,)�?(�p^�SP� �#AY� !��bs�ADc ���EX� IO?���w2�b%JQbA�P�a~�fWR���)�D��v��,�F�RIE�T�U/ M��$TpTOOL[vM�YH� �LENG�TH_VT�DFI�ˡ�s�= 9 �yU�	@V_{��p�R�GI�cWAITI�N1��uX� �z�vG2�gG1�a ?��rb�P<PVr�O_�" C@�@tqܠѐ_��c�%��ATC��r!�]��qGÀ�#AZ @�� ��i 2L��h��!���!D���� �d[�X �"MXC kP9����h����d�c%G�Wh��""��DEAD��K�D/ELAY8 T�!2��F��!  x� 3!Z��q�y1#xpU2{2��3{3#z v�͑$y���,��`��L�`��$V� �rV�u�V3�su�=�� \ � �_�e�uc�L��Y�B��T�QR����Q���s";�$`��PR.P�����S)�.���d��] 2���˃k�[]`2�k�\;!{ �0���p�
��̂S��^� �@�R2��7 n��UNN��AX��;�A�pLq�2T�T3HIm�2LI= �FEREN��Q�IF�PsT�Iw��,��(�G1����+�ĹA4�q?�ܶ_JX0��P�1@�p�TJ_� �T R#% �2BD��r�C�C)�B�Uy �wq&Q�5�Q��#IN�W�p��$TBC[_P�pCM�#DW�2LDR� ��Z1����@��iCLASWIT��C0ATA��`�"��D# �$VA�LU��O���Np_ �a����  2`� �SC��b	�� �$ITP_�d�BU$�TOT�K�$�� ;�JOGL�Ip�	A_PJ��O�e��c�0AX�P�K�`aMIRW�w�!�ML䂘�AP�!��E�A�2�QSYS�шVP�G��BRK5�3NuCK�I<�  �Ҁ�#��&���B$ӑ�B#SO�A$Ӈ�N+�#�6�!@F1��,FS?PD_OVRwp@����LDf�i�ORt���Au�F��u�T�OVW�SF��� ��bF��R|�%���eq>��CHDLYq�q2e�@T�W� eD�W��RO�7�c�3 # @p �0�pE���10�1I@��Y3WD�!� ��7��b��Q���F!�AF4A��)�y��BB�2�P�%�"Q�ˤV)4��Ӧ�3P���A�M��)��  ?�_�M��M@{L�T$�CAJ�[BóT$H�BK#2f�!s2uI@r��PAi
��z	��%�K�DVC_DB�3�Sp�� ?W�1�
?�3$�E�A�`����f�Us��{l@AB �r�C=T����Z1T��_AUX��SUB�CPU2bSn2S�c��j ������F�LA�A�HW_C v��M��\�A�@���$UNIT�| �ATTRI�М"bCYC�@^C�A;��FLTR_�2_FI��TAR�T��p@B�bi�L�Pm�nACH_SCeT!cF�0�F_,��"*FS`!*2 "C�H0t)�!�D�%RS�D4��jyA� _T���PRO'��n�E#MPI�4���T�"�� �" �B5�PG~��RAILAC��2M�LO�wsC�5_r�QF�RF?P�R� �1 ��1C�� 	>�FUsNC���RIN~�0z�W0�4m�RA�0:b� c �3�@_�3W3ARճR BL�BF�'DA K!#HHDA`��1aH'C ELDW Y�%��C<� A�Q�C�TI���E�a@�$�πRIA���CAF�P��`�A7��E���8�zU��OI ��D�F_}p:�PD�BL��Q�qA%�HRDY�dO�Pt��Psi@(UMULSE}p�ө*)�C0Jq�J�����FAN`MLV���QWRN�UQ`D�,`i���22�QST�O���_���AU�D�����`O_SBR�eH�j���1�4cMPINF>�p!GdARcREG��cNV"P�c��DAhp��FL��$M Y����W? @��X�e�CM��N��Y�3N�ON���\� q���a��c �vAq$��$Z�q�����d$ ���EG��2�Y�4qcAR6�J�527K�CuM@��AXE>�R�OB;�A�;�g���_�}�SY�nq�еvS�wWRI%�Gv��STR:�C �Ѐ�E���Pt8K��Q���B�pK��9}3+ O�TOba���@AR�Y;�=�w1+��l�FYI�Ђ�$b�KQ�[�]��_�sK��B�3�0��XYZp�R�����OFFS�R\���x�A�B9Ђ�2�����0�F�I`���\�Q��2�S�_Jf���~���$�P��3�$�US��B3�fRk�CLQ ��DUg"�53ҡ.�2TUR�`X�C���K�BbX�pY S�FL����ZAp���3�J�a� 1c��Kc�M�Ԓ��6����{�ORQ6H��3Y�6�5��ѰP�Ar���8F�ya��OVE��^�M� бs��s��r ���P���Q������ �0�!�@_������� б������1�s1�̣�H�ERe� A	�2E�%����3o�A������52I�hAehAAX(���hA��>1_�ɵ J1չtQչJ�Ժ�0Ժ i�ԺWpԺ�Ժ-�Ժ1��ԶTPѹTP�TP �TP�TP�TP!�TP 1�TPA�TPQ�n�b�@ �R��DEBU��$�1�SB2"�h�A!Bh7f�ሣV[ � 
=��I�e�� qכ�q�J�q׉1q�i� q�Wqq��q�-��Dp���B��LAB��8S���GROT S��\D B_(1V��t ���`�N�T�J�aV�AND��d�E��g�a�� D�a�p`��*A��G ��NT�`���VEL.1���0f1��2��NA����rC�!��c�Wsb���ME�SERVE��#pe $���0�7!_�PO������7�f� N��"p�f�`$��TRQ"��
��r��g���B�2f���@c0_ �h l�0�u&ER	R�;"IY �����'TOQ� �LrpӴ(�r0Ga�%r�x"��`��REj@ i� ,]����g�R�AI 2h d�f����� j�p$��-2
Pò ��OC*A��k � ��COUNT~�q NK�S�~sl� �Q�MS�f��ELAYt'�VA ����@���Q�A �1	mfCS�`>�EKI#Xq(VqVUSVSڡ�HFX��Y�ZV�NU�V�W�HPK2ű�C� p'p'~'�'��Q�SFI4�1IG�@DO< <��M!���K#��g��2�m� ��,�c	$NJ0 `��7�SFJ��7�L�FZN_CFG��n� �`}d�`pcFL\�Q���� n0�#so{ �b�MIN_�R�I��0����,0<5FA�@��F@3X�pb;<9�H�}qb�$NEz�qP�R4�SG�@�GOUU�p 8��`arO�S���0�Bg$CU�P�PAj��DLhv��1THK�CN��q �b�Gf�`HK3��AG2KCUN��G0GC�8IPGCSEV�BDpESK�P@�aJ�Cg_RQ�R�7RP�2�r\ $ASES��T���@I��pc:��DTRGQ�BOBSrAK��`��F���GCL�@IC��CX��$Xm�X�{�@0_D��?SF��=TPL2>S�@:UQ1CXuPQW1\Y1iYQ2CX�PQW2\Y2iY/pTDOW�[0�S#_O�crR�ACp�4�Q�WA�2MP�a�Gs (��� �`1��-c�`6g3�dST�U�at `,�P�0_SCHX�K�W7ELDw�ESlS|b�MW`:S6�EW�UR�=�@%�_!����� L�L���RfA�1u� ��� U tޭ2GDTP^q v <�0�0�����:n�AX�\�{��u����4D�bw � ��/W���icuWTCW`�4��zu3�u��H�GUNat$��3S�s ���u���ụWD�*u�1WT7vx��d�`yv�bp�3w d���q�dy[��p_�,j7�@b�"HC�$�z��@CHG_PHAS��$��$�`�P���H��  �l��d�C�� @��AV�m`L$P7�$WAITT��T�pru`�A��PWU0A���B���LOL���Ƀ2�p�C�RIGG�EREW1$KE�EPa�?�$SVqO�0���CAL�c���A�R����TT<��POWR��!L�߁LO#RpO��CTL� ���n@���IOyp_AL�1�EPOY��{ � $Z�%ӑZ�b�P��	ᡲ4�������_BY�">�Z�S�Hn�$AUTOGREFc"6בCs����VIRTUAL�\6H_6��avMKUL��GA�1H�a~�#| 5�wB_BE�RSR$�#7$	��*�10�2�3�4��5�6�7�8�0�RO�6גOmN�2$�1ABp�1��N�IN� ڐ�����2�S�� ��_�PUQ�!���0esNS�$��a1�"���S�PFWD_KARH������R���O`;ON_SQUE��x��D�"Y�3C�0PI��Q�ΣEX��ɱA��o@Mmє�{�́817STY��SOP$��DI�AM�JuD�IKNI  M|�˂NP��Ł�E�0�eKEYSWI��i��!��e��HE� BEATM_S�`M����K�6�Eؤ�0�F���S��D/O_HO `S�2��EF�r�� 2��Bή*�8EIO��S���P_IOCM�qm����2ϣ�A }# Dd`��0U��Z��`-�PO��$FwORC��WAR�Q�QPͥ� V�~ @�d`FUNC�CćPAR��b�@cf�Mbe�}4�S_R�S� �O$�LG�R��UiNΑ���ED`��0C LCLp���l ���ANC�ELp���I��ؑD�RY�����WET �%��������@���81ZON1��^�V�U2f�2V�3f�3V�U4f�4V�5f�5���_SW������PcUR_ 	��SEO 0ؐ/.�EQ��Q@.��6=ulY�ѱB|���RS��O��@���U�DEF e�������������4���T�6��6�7�7�8*�8�9�9��.f�Ee�#*�� 0#*��L#*��h#* ���#*{�#*��# *��#*��#*��3��GI_BCK |��`%<$5��18L5$5��E18l5d6'�6��!O딚�7�6T}Ұ6`�3�8�7�8SV�tI�5B��H_R)��#H�5CLR_XF��?L>FY\��bI�5X1�L�5INeAL�6 �E�G`��G�L���G�L ��W�L��$W�L��DW�5MAJ)p'�dV^W �CmW�C^V�@jY�S^V ��x�mV�T�Z���Z��ƺZBYmFe�WT_aN���W$c�5NO?� p�>i�5��Ҁ;`g�5ROBH�D�g�5 6���5�e�5��g�l �F�fV$�f-VD �fMVd�f{`w�l� �w�l��w�l��w�l �F+��3�iY��w��PL)f"��f(@�:� �F>)@�VZ)@�-Vv) @�MV�)@�iv�)@��v �)@��v�)@��v9@�8�F9$@CKPC�W��R�EQ:�b�z�R�FA��b���R�L0B����R��hADb�ЕȚDA���R���^�����8N�w�����/0���� 9B�0/0G�ROU��LAST�_BIT��v�r0E�RFa�EG�^�_T��>���IN��H����� I����O��H'�?��V��ݰSeC�M��ߡE_WID�T�M�N�SIZ �`#`[ቢ��ϡ��TPҪ����� �FIGt�����&@L����r0��f����f�3p�4v�~�TO��  	�2��6�AIR��F�}��X̳�2��EF��P��:���TOG��"��CC���G����SPX\�&���$ŋ�#�T��#�5 �6 �7 �8 �9 �l���}��� ������`���m��� z��Ň��Ŕ���0`����֋�֙�� `��m��z�և��Ɣ�O��Eb�� � �ѧ� � ���PSCF�G�� � $r��D����HAN������_CTR�$�IS|�#�T�IE6��PD��SA�ڴ��VO_TYPE %��	俠B'��Ѐ��x�9���F��F� �4�SMB_H�DD�� � ���BLOB   � �SN%�A�S��� 0 $ADDRES���$�$VAR�_NAԱ%$M���PLYiё㠠A��� � � _$TIME��$��;_I��	$������⿡CI��FR�IF��N0SION���U��$�IN�FO����BUS_GADR�I�D�PHd�$CMD�`DIAMN��$zA�A��$DUMMY1�������$R�A�PCi�o0��� @� ���y�Q����URy�NC���8�������SWi@��� L ���ЏGRP1��� 2*#3#4#5#J�~�pT � ���}S��LESTEz�|���$SGLp�TASK'� &�/�����q ST�MT#�PSEG�#��BWDpSHsOW���BAN� TPOF�������0��a��SVuC��GV�� ���$PCz@e`��	�$FBiB.SPCT�. DRV��� �$���A00'�+�p1�v2v3v4v5�v6v7v8v9�vAv7�yCvDv&�yFv:(��1���:(�1�1��1�1�1�1��1)1)1)1�+)18)2u2�2��2�2�2�2��2�2�2�2��2)2)2)2�+)28)3u3�3��3�3�3�3��3�3�3�3��3)3)3)3�+)38)4u4�4��4�4�4�4��4�4�4�4��4)4)4)4�+)48)5u5�5��5�5�5�5��5�5�5�5��5)5)5)5�+)58)6u6�6��6�6�6�6��6�6�6�6��6)6)6)6�+)68)7u7�7��7�7�7�7��7�7�7�7��7)7)7)7�+)78$$\PR�����a ����p��� 
z�V?�`� x $TOR����D�ะH�"�=�El��-�Q_��RE0F/�AX��ݰN�SE��CARTY� v�_�U� ���YSLO~��� � �� G�0���9�q���oVALU��OP?����R�F��ID_ILC��H��I��$FI %�8����$��q⚃SAV�`� h�c�[�L�CK5�p��y�D_CPU��������4:�L�T��TE�����R � � #PW����LGᝠ�Re�� ���RUNB��G������W� �7���7���H��X��0���T2@�_LI����  $eJ��O%��TP-��DIRq�SPD6y����EN���������k��TBC�2b� ���E�NB��I��y�FT�Mo��}�$TDC�����M@����TH��.�9�:�!R�:����E��\�p)�\���͡_AC1�� �X -$��LEN����)���EL_RATIC�$��W_U��14��$�2ηMO����|����ERTIA]�`0���"����DEž;�LACEML�CiC�_�V��MA��p�T�*�T�TCV[�|�*�TRQ{̜Œ��N�*���*�*�J_$0�2M���J�`R��*���2��`����;�JK2�VKc�D�)�Dњ�9бJ\�H�JJP�JJX�AALH�~�PӐ~�x֦�|�59���N1�̯�n�X�]� I��� W YΠCF��7� `�GR��V�(� E�:N�C��v�?REQUIRG�9��EBU���$T�3�@ᄰ*�͡���Ӥ� \ ��A�PPR6�CL]�
u$��N}�CLO�����S$����
͡P�ARA{�� � M�k���Q���_MG����Cbd���0�h���BRK��N�OLD��� RTM!Ox�3� ���Jx�2�P��6�P�6�X�6���(6���6�6m�7m�~�R_P��Ӥ�G� 3⮲c���<)���PATH����@��������E��r�SCA��6�~���IN��UC���F -CPUMOYаH�1�V�b�q
)�q
���q PAYLOA�.�J2L�pR_A	N��L됼	��	����R_F2LS3HRV��LO�E��SSACRL�_y�C6?�Q�H��]�$H��dF�LEX��E͠JѦ� Pj����[��m�W�_���� :����*��$��`R�*���ÿռF1! [%o'�����,�>��"EH�Z�l�~ϐϢ� ������v8�4����2Ԁ� �8����!$�T�t1X\�}10��$8 ;�DE8G�Y�k�}Ё� ��x՜ե߷�����Ԑ��ԛ �ݠ����|��pAT�&2���CEL� ȡZS9�JE��@�JE�CTR�?�!TN�VV*�H�AND_VB]������� $�0Fi2��&�߃SWV��ʣ��� $$M� ��7��h�l90
e[�5fA�� ���Ri��A��Հ�A��A*�]`�뢐�D*�D*�P
 G��iCST��a��aN-�DY�{���>dee�  ���!��2��45 @1�Pu�~��������������Jҥ�c �P��� �!x�u���ASYM_�3��a�6:_X�+K ^H�J�@�Xhz���J��h��
�߉�	�$_V�I�S&���7�V_�UN��%�L�mC�J 3�d��ud�h�u� ��'��:h�I[��%Cqy���TC�PPIR���  䰦*0P(Џ�CDELAYnA��D���G� X��7�@NȠq@D� ��l�|а��d��!�0MPeRP�ROG_t��PYP�Eȡ�_T� �7���-�SE.�S���BಠRVWARNI8{p��OTF�!��f*�_TU�MAk��ޤC�VߠABCF�IL FQ��DB��Ң��
laMPs�I�Z��l`T�X��ARExr���������REչ�~�������_HIST_BU�_ � ,�0P9PQWPR���t��uCI�DT� �P�7��PEARTBE��SETPP��.�gARGk�*�FL��\sţ�STR��������ŏ���������(�OUTO�� p@�m�Ti�E����ܢF�ID�@�U�# 10�F j�ieL�ҤA!dX��pH�o���Rtt��Ii�$DOi�r�P�t�S� }@
lbIO�A&�H��Љ �t���� fP�P� �ߨ � �QMEJ�!��R/�t�T��EP"��j��D�����1�%�T̀�A� $DUMMY}1��$PS_� �RFH   ��l�4�FLA��Ն�$�GLB_T `����@��2��P� �Q�ѩT�Y@X��ST�!P�SB��AM21_�Vz2T$SV_E�R� O������CLĻ���A� b�m�GLv.�EWO�� 4V��&�$=�$ZnBWJ�1�up�SA��O��,�U0�� ��N�d�Ҁ$GI�P�}$0� �8*�c�O�� LV������}$F��E��N�I�� N�#F��� T�ANC�"B�J��R�Ra ��P$J�OINT'A�@�*�MV�O��"���E���!$PS+R)�$QO�_��  � U�!�?�PLOCK_�FO�Q�BGL�V�SGL~T��_sXM�=EMP �z2:�� ��i $U�/�O 3�Pc������Pn ����CqE�@���  $K���)0M��TPDRA83���VECD�� IU���HE�p TOOLO#<VvN$REIS3�2\6�qr�CHV�{P��z�N"�[�3����SI�  @�$RAIL_BO�XE'APROB�O�?���HOW�i��ROLM t���A��Q�w n�pO_FP!P�HTML5��S��JU�P+R�,�vO���	&�R!OCO��N	SLO '�N�Ĳ tP��S°aQ:Qi �"POr!��IP�N�0R��v'��I gCOR�DEDn {Ph ��X	T� 3)���a�O��� D ��OB�adSn 71U�Р�2��fQSYS1AsDR���TCH$`� ����Au_�s4�AFQ��PV�WVA�� �� 0�����V_�RT�q$EDI}T�6VSHWRQ�@V�0IS��B�I�ND��{��4bBG�D���@���3�KE=�O�*�FJM�P#0L��W�TRWACE���0��I� SeRC�PNExEfQ�WTICKFbY�Mڡ�rICHN��� @0fAש_qG֧�4�STY�{�LO����IB�B��P�� 
�%$Ԙ1��=�Sx�!�$Z�F �ս��P�<�צSQU��ԳLyO�%�TERC��ԱD�S��� ����t��/ ���	T3eO�	�װl�H����hᖠCt�<�R��UTPUQ��Ug_DO��r0XS! �K��AXI`#��URް!���$T��@16Y�FREQY_3C2ETDbPw�0�\�F�PA�,q1�\�9�2��� SR�t�l�P��:�SrW!@Jq����iq�nV���fNr�hAxp�gC�|A�pAV��u�b�6z�a6xD0~DB~DHT}�5yC�C}CT}�������τ wPS}C�� � h #DSh�[��X0�c��_� d���pDX�AD�DRESFB�0S�HIFPÿ _2C�HB0-1I������TU��I�a �>i"CUSTOed��VSI�ҽ��~b���`
�

 48���T�о \���(A�\�ӌ�QB��Cus��Rhb⊚&���T�XSCREE2�z��QTINA"���c���m�EaE��0� TXA𧥧������aB2b���0RR�OR_��d�������UEzT���\1z�S�#�C1RSM�@gU`� nP���t�S_]�:��S*�=�X��SEaCxc��� 2�^�UE�c´��}�>�PGMTN_����!`��!W!E@BBL�_�WB��� ��\�ڢOW��LE�u�����RIG�H��BRD�k�C'KGRB�"�T� !�>�WIDTH��0����F�U�I EY, ��� Ad�����B��QBACK�At╵����FO�!��LA-B�a?(��ID g�$UR�հAC�m���HБ � o8 $�T_A������R�0i�c�Hd���O|���ƭ@I��U�F�Rw��LUMF�(fe�E�RVO�l�P��u����y`GEٲ��c`L�"@LP��nbEkP�q)��������p���5��6��7��8 ��iR�S�P��$�Z�p�aScP�m�U{SR0�� <��b��U�򸃉�FO��.��PRI�am��Qޗ�TRIP�m��UNDOMDɂ��'P�Щ����q��B`<P ��\b��QG PT ��q����OS���R H`֒��B ��9�K� R�*��D���U�� ���3�E�S���KU��OSFF� �0�(�[�=O�� 2� ��Z��� GU=1P���U"���q�炱SUB��B RE_EXeEM0V�A��WO�a� �z���bWQA�0b�%���a��V_DBD�\�SRT,���ϭB�� �SOR���RAUD�`��T��[Gr�_�0�ND� |�`[HOW�N� z4$SRC�ᐷ %PD� ���bM�PFI�D�qD`ESP�Q�R{�Tu×q��bW���0��� `��2�z4�QIPCOMP�1$�@��_ `��!�N�CT4��2�@2�b�DCS��Pc"�45�C3OMs�qPZG�S@�Q�E�Q_�Z��ᬵG�VT�~�
��Y0Z���b]P�=Q΃SB;SU���" _#0MA3|��0gDICv�AY�.�RPEE0�Tڱ�Q#VR�00���p���Z��S�� n���^�L��+��0�� �� ӣ�SH�ADOW� h�!!_�UNSCA�1.#OyW�" DGDEv��LEGAC�ȇ ��VC�`Cs��� �B<1?S� �PAR���,GQû�C��^�%DRIV�VOa&C�!@���6�?MY_UBYBԖ$ 	V*�?U�HP{�@7DG�1_7 �D=2L�[�BM�$q@DE�Y�CEXǠ��M�U=@XT�2/�USAA/`��_Ry�ZR���zp�[QG2�PAC3IN�A0PRG�4��2���2P��2b��R!E�y�*���s#�2N~P� ��x G� !PF�@��t#R�~PA�}�?�ϑc��	��aRETSW�0_IA�1:�3�POXѢk�A��B�bE�PU��@� "�t#HKt��<��J��a8�@���CEAN�I2�����E��t"MRCV� �� ���ORG`���	R��CRREFƧ;V"VQx@ ��rc`@g�ZqQ/ZqQ@[�U"V�O_���J�X�K	pS0К�#��t"��� �7�$�VB0h�s��%�OU����# �+E�q2�ա�d�&�����`D��q]a�e�ULv���E CO���s0p`NT@�dN@�e'��fOѽc|`L@��eG�e'��gO��wVIA1�� ���HD����$JO�.�Ƣ�$Z_�UP��Z_LOWLuq{c �����$EPpa���<q qW�^�s�^��@�#���� 5D�PA�O� D�CACH}3LOeQ�t�qt0�y�Z�� C�Iv�Fĵ�T��k$H	O�����p��#�O�J�,gc��c���0d VPB����_'SIZ}3��Z{���Lq��N�5�MPF�AI�Gm�pA9D�MRE/d����GP�i0 �A�SYNBUFR�TDD�P���5�OL�E_2D_��l�WHP�� � Ub3�pQ�@�4�ECCUHVE�M�0�u���VIRAC�d�L��P�_�����Ю�4AG`�R�v1XYZ\�D�v1W@FA$�cQ#���ѐTy ��IM
�c��Z��GRABB'�S�@�LER�0Ce`�Fc_D?0�q�50��H@���
�uz��p ��LASP�IQ�qw_GE�u� ��@Ւf��T  y!F P��5I,�B�� ?BG_LEVű�!�PK�0��,gGI��N���B���p$��p޻��qS��vIN�� L!�t�"���z�f A�y�D��DEp�' �Y4nE3p�� ���n�AѺ�G�O�9h�D���p!��T�Un��� $=�IT����в�5,��VS9F{ �s�  �І+̽av0UR�B<ASM������ADJ�t��pZD��� D5�mqALVp����lrPERI��$�MSG_Qd�$@��ƅh�N��r���������up��^��XS.��� x��M���dmqP�P��<RSM�нBlrLNTK��M�,���ՅC�pAC�&%`�����"n" �7XVR���ݢ���T_�ز�ZABCԤ�'B0���ZP
�q	�ACTV�S~p � � c$Y���Y�IV߱�^�IO�"��Y��I�Tl#�2DV& 
H�1p�
0݁��PS �^�8���^�LST�^��pd`��_S�g�SGT�� CH���� L�����OG� �s[ �P��GNA�\����^�� _FU�NVP^�`��ZIPf��럲h'$L��ZP�ZMPCF4��£���&����!7LNKB
C���~5�� $W���@��CMCM�0C��Cy��GTPX� �$JD ��,%Ǡ1Ǡ0.P5T*]UX/���UXE�1}/� t�6t��	�� F�TF�a�IQ�=Zy�� ����q �YupD~� W� 8�@R �U*!$HEIGH�3Ƒ�?(x`~�YQT�I�d� � ��FQN�$B|`%p��"rSHIF$��R�V�F��ZR�%�C 3p�d���2��������D���CE��V%��SPH�ER�  � ,�x`*@R����T�HRSHD  ��� F@ ��]!M!QZ_�ED��  ����e)TT��q 2$"�'� �#
�/�/6�/ 
�!_A�Q��T��#e%�"M�@<H�z#  �*�0؈�/m!UAy�PL�5?i$NO�pCK ?�+����$�8�? �?�?�?�?�?�?OO ,O>OPObOtO�O�O�I m1Ԃ��6�'m04��SP   �-x�$_T�$ODh�8��5A:OFF��/�8��Z?IWDISW_HS�=� ARK6W�)OPEN)���z"�!�&�)Q��_IO6W bh"�RW��`%�*�%$*on�S"q ��%N�"��If�#�!���  � ���$d`	Qlf 	 ���F2cb�F�C��*P��DSBL�  �%g!h]��o�LO:�NTl�fZ$C�0f!A HR��SIM_D�Wd�"Da(*P'�SL ��+}$]d]�edFT'�_P��w_jv��7Vde%lt��3~O�� ����t����AM2c� 1�xw��s\fp vgR�d�v��������� Џ����*�<�N��`�r���������̟2 H����'�9�K�]�o������"����ϯ ����)�;�M�_� q���������˿ݿ� ��%�7�I�[�m�� �ϣϵ���������� !�3�E�W�i�{ߍߟ� ������������/� A�S�e�w�������@<������/� A�S�e�w��������� ��vfS�����p���"PI[m� ������! 3EW&8��� ����////A/ S/e/w/�/�/j|�/ �/�/??+?=?O?a? s?�?�?�?�?�?�?�>i�/��	Q�O 0MbtB@OOaMEO�O �GMM{C�OO�O�O�Ae`vg___1_ O_U_s_�_@8p�_�\���E	`_�_o<o�Q:�oq=o0Ooaoso|@Bp�i�G��p�c1rp�RM��@�$�bW�  �Z�p�~q�h�O�O &8#\G��}G� ������ �2� D�V�h�z������� ԏ���
��ӟ@�R� d�v���������П� �����*�<�N�`�r� ��������̯ޯ�� �&�8�J�\�n����� ����ȿڿ����"� 4�F�X�j�|ώϠϲ� ����������0�B� T�f�xߊߜ߮����� ������,���P�b� t����������� ��vo�e��T�x� �/������������ ,>Pbt�� ������( :L^p���� ��� /�$/6/H/ Z/l/~/�/�/�/�/�/ �/�/? ?2?D?�Oe /O�?sO�?gO�?�?�O [?q.OORO	_�_}_ O�O�O�O�O�O�__ �_�_N_`_r_)o;o�_x�_�_�dA�  �Y BOo>L�i1o�o�_jo Uo�oyo�o�o�o�od���$PARAM_�GROUP 1�!�!�|� �ERj5 �5R#q @D��  7q?�=s#q?hd�?q?�C�PEzYs����o  ;�	l�Or	 �`oL �p�@`�A`�pX0&;��p� ��rP�H�mH����r�/H�cH,���l=�oy?J��QB�P��)��Wq6��s�4  �Z@p�=�ôQ��Y��?�Q�c��cBR�B��Ϯ?�Q	�;��2Ǐ͂Pq��#oAo�v�  �j�K#��  ?�  �/��o�M��u	'� �� k�I� ��  ��U�v=���͏����r@������~)q�R�)r�����wN4�9�  S'O�PCx�B��A�Up��B��k�'��_�q�B� ��{D/�y��3p~�| �}��4����]Α�?�D `u<�9�$�]�H����}�O� �� Ơ��[`{�����3  ,�d�:fu=���@0߱?�ff0�?����� 4P4��F��q8d�\�j�>���Kq�z=	_  �����P"��ü��q�s�t�>L��q��hQ;��~�;DA� �g;�-�<��ް�^O�&���Or)s���P?f7ff?ΐ?&I��t�@���[�A
�g�ٳ�D�Pt�y?u ��=w��-׃t����� ��;�&�_�J��� ������������� �߮��m����|��� ����������3 WB{f��tj 0��T��ASe,w�A�y�Hϟ�R�B�<���0�/h��QA�A$�YT+C(���5}/�3
���,?��@I�ܦ//�/�/w�č��Sâ�܄��pD�9p;���
� +�� ���/�rD\Y�C��s3C��B�33BZ�P��h�� ���� A�333����Ù?��9�3�ٙ���_��Bm��A�33�?���0;�0nffBd}� ���[�<PL����L��K3�ÜIĮIK��G�d�� A��3,L�4L��ʖIb� I-ߞ�G��:O���4LA�L�?��I���Ir�H#Ο�O�O�H�71�O�O�O�O{qA{�?_0&_/_h_S_��Sv__  F�d��_�_ J	)9��_�_J	��o [_4oo0<?Foojo �o�o�o�o�o�o�o! E0B{f��~ k1����b" ����?����_O��?���n�y��1����B8�ޏɏL�Z�_��� L����KI�6�A�z�e���0����ԟ��G될���D_�K����J�5��n�Y���}�����Cf�Ưǯ����2(�13gf������G������7�I�̱q3\�o�5�3|����5��L�|3z�	���ͼD���E�w3��� �'��K�9�o�]̘%%P�P�Μ!��� ��� ���$��H�3��l�W�:��~ߢ�1�E��e�������� 6��ϯi�W��{��p��������<+J����� :~ �����W�E�{�i������  2�0�bGC�\(��B�I @!�KC�50I �0@P/ '9K]o��#-�����a4P���$�!�$�0���s$r!�+
  �\n����� ���/"/4/F/�:��%��H稤�$��氖��! @D���!?��! � `?d1����%�
�,�;�	l�"��0 9��,�� d<�0aG��)?d/��W? i<ء��?�9�?�? ��?�?
O�$P�+O�9H�7�����  ��{O�H�?�O��O�O =0�O[@��1��_'V��&ܠ�A_S[�"��{_�'8�_�\�0A��>��_�n_�_����<?o�8BYo �oe��EC���_�o�_�o�o|�o�o �c �1$w � ��:JbA$6*H?q�"�lL^�o Q���{���8�0��z>3���!ߚ�.o�>L 2Br�1T��u����#�"l`?fff?�?&���oŏ �������6�%���( ����$��S�>�w�b� �������������� +��O�:�s���� l�ͯh��ܯ� �9� $�6�o�Z���~����� ۿƿ`O�Կ5ϐ�V� ��}��ϳ�����v� ���Ϙ�1��U�@�y�
d�����D��Ѳ� q�����j��/��!�� E�0�B�{�f����� ���������A�,� e�P���t��������� ����+O:s �p������  K6oZ� ~�����/� 5/ /Y/D/}/h/z/�/ �/�/�/�/�/?
?C? U?@?y?d?�?�?�?�? �?�?�?OO?O*OcO NO�OrO�O�O�O�O�O _�O)__M_8_J_�_ n_�_�_�_�_�_�_o@%ooIo4omo��(������o�k�o�o �o�o�o	�o- cQ�u����|J��Pg�P� ��� `o1��h6�`�K���o� ����̏����ۏ�&� �J�5�n�Y���9��� ş�ΟП���<� *�`�N���r�������pޯ̯��  2�� 6�H�Z�l�~�������ƿؿ�%�
��.π@�R�b��Ո��ϖ�
 �ϵ�������� ��/�A�S�e�w߉��߭��r�����}���$PARAM�_MENU ?���� � DEFP�ULSE��	W�AITTMOUT�
�RCV� �SHELL_W�RK.$CUR_oSTYL�I��OPTA�`�TB�t�n�CD�R_DE�CSN�SGT�IPCMP.$E�QNUM���G�UN����PR�INDEX�M�ISC[2].$�HPD_TRQ[�1]�����1.$SETU����u=� 7�I�[�����������������SSREL?_ID  �������USE_PR_OG %��%��E��CCR!�����X_HOST !��!]�R
AT�d�}��|�Q_TIME��m��GDEB�UG ����GINP_FLMSK�JTRYJPGA�w :�ωCH�XITYPE��������/8/3/E/ W/�/{/�/�/�/�/�/ �/???/?X?S?e? w?�?�?�?�?�?�?�? O0O+O=OOOxOsO�O��O�OLWORD �?	��
 	�X�}�{�AL�!�	JO���CT�E� {��ICOLPyżHG_�LQ��՜}��md/TR�ACECTL 1�����	 ��� �r�� ����#�r� r���_�Z��VDT Q���`�PD � �K�� `
�dddd d��b��b b�bFa��gbt��b7bHd�d�^a� 4�d5�bG� �d���b�dU�d�d �d6�dU7�d8�d9�b��dU��d��d��d��dU��f:�d;�d<�d�=�o�o�o >�d?�d@�ds��o	~Db �`Lb�`Tb�`\bI[��ldb�`|b�`�b�`I��� J�d��b@?P�b���b���bO�$�	� � �bQ�dx"�bS5�G�Y� !��bU�dV�dW������� �bY�dZ�d[��d\�d�b^�d_��d`bJkc��tcJ �Q���Q���Q���QJ������cJd�JS����b���b��!Teo��"��#�������da�db����џ����$cJ &]�'J]�(]�)�_�*]��+=��bc�ddb^�c�^sd^s�^{�^���^��^��^��^*d^d^#b9�K���l,�d-�d.�d/X���	� 0�d1�d%2�d3dd�Ksft�UK{�K��K��K��YK��a���d��d��U�4�U�<�U�/�[�%Yļ�U�Ģ U�̢U�ԢU��U���TU�������kc��tb��t���|� ���������������� ��b��b��$b��,b ��4b��<b���� ���������*������Y����������U��cE�d��d����U��,s�3t�;t�Ct�t��t�s��{�󢃄���l��s��{�����S�� gY�hYĂ�YĉYĊYċYď�YĐYđYĕYė�YĢYģY�D�U���YĲYĳYĶYķ�YĽY��Y��Y��RY���� ��Y��Y�)�)�[�����r������� o�[�����`�d[c�[sd[�s�[{�[��[��[*��[��[[�[��$cU[+d[3d[;d[W� ��`���h���|�����T���[�[�[�T��[ä[ˤ[ӣ���[�[+s��4sU�7��G��O��W�U�_��g��o��w�U��ׇ�׏�ח�w� m�� !P|�$t�&��AP;��8|�׃����kc}tb}t�} |�}<�}��}��} ��}\�}bim}$b },b}<b}8�,�P>�P�b�������U���W�ô�{�1�a����Q���-�,�/��jb�/���+a??+?=7��`�GԼOԼWԼ�_ԼgԼoԼwԼ*Լ�Լ��A0X�G��1P�4 987:�9X1�Ӻ2�5 �7A0t���!O3OEOWO iO{O�O�O�O�O�O�O �O__/_A_S_e_w_ �_�_�_�_�_�_�_o o+o=oOoaoso�o�o �o�o�o�o�o' 9K]o���� �����#�5�G� Y�k�}�������ŉ�)�/�/������-�?� Q�c�u���������ϟ ����)�;�M�_� q���������˯ݯ� ��%�7�I�[�m�� ������ǿٿ���� !�3�E�W�i�{ύϟ� ������������/� A�S�e�w߉ߛ߭߿� ��������+�=�O� a�s��������� ����)!�3�E�W�i� {��������������� /ASew� ������ +=Oas��� ����//'/9/ K/]/o/�/�/�/�/�/ �/�/�/?#?5?G?Y? k?}?�?�?�?�?�?�? �?OO1OCOUOgOyO �O�O�O�O�O�O�O	_ _-_?_�O_u_�_�_ �_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o �o�o�o%7I [m����� ���!�3�E�W�i� {�������ÏՏ��� ��/�A�S�e�w��� ������џ����� +�=�O�a�s������� ��ͯ߯���'�9� K�]�o���W_����ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g�y� �ߝ߯���������	� �-�?�Q�c�u��� �����������)� ;�M�_�q��������� ������%7I [m����� ��!3EWi {�������� ////A/S/e/w/�/ �/�/�/�/�/�/?? +?=?O?a?s?�?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O �O�O�O_#_5_G_Y_ k_}_�_�_�_�_�_�_ �_oo1oCoUogoyo �o�o�o�o�o�o�o	 -?Qcu�� �������� ;�M�_�q��������� ˏݏ���%�7�I� [�m��������ǟٟ ����!�3�E�W�i� {�������ïկ��� ��/�A�S�e�w��� ������ѿ����� +�=�O�a�sυϗϩ� ����������'�9� K�]�o߁ߓߥ߷��� �������#�5�G�Y���$PGTRACELEN  \��  ���\��q�_UP ������̨�����q�_C�FG ��,��� ���[�\�A�����������������DEFSP/D ��&�����q�H_CON?FIG ���W \�\�dg�MȀ� &�j�P������\��q�IN~��TRL ����8���PEL��V������\��q�LID�����	��LLB 1�V� ���B�v�B4F�� ���_Y���� <o< %�?�� �������& >\BTv�����r/// D/�=/z/m//�/���GRP 1+��\�D/�����33[�ALQ��IK�HU� �I3�@Av�D	����k���9-9f�f�� �/�FI>´�3b?K;B�0 �1�?t?�?�?�?�?[��C$ 'C*���O;OMN7O <C�rARO�ONO�O�O�O �O�OjO�O-_�O=_c_DN_0z�S�_\�
x_ �_h_�_�_�_o�_7o "o[oFoojo|o�o�o��o�o�oz![�
�V7.10bet�a1�� ?��?}?�-@(���D/g�D���D�vfD+{R-6qET� ^q�D��[q�pfE����E5#�C�� 1C1GpFt� ������A�p���2EJ�X*�׮�vD��A<>���B�F '���F l0���BO�33�Z��Z?�:��X����� �o�?�o�6j�|�f���$���.yg��";2e�Ə$������-����7p@�!�p�r�� �B�BQ{�m�BHT����\�\���6��������ps�ΗD0 �B��<V�E�x�z�<��r6�D�M���C�ԼB���
�X�R�i���A�4�j�£�r�2�f���������r��������?+?=4 B�S��w�b��� ������������� =�(�a�L�qϗςϻ� ���������'��$� ]�H߁ߘ_�߷�f��� �������5� �Y�D� }�h����������x�"HsF@ 6� 2�F�X�v�������� ����v��!3J� W��{fx������@1u0�R�4� X�m��������2K���0���x�x>�: /
//Z� 2&g/]/o/��/�/�*ޡ�$PL�ID_KNOW_�M  5��1�$SV �2%�  K����6?H?Z?�~?�i?{?�?��!��#M_?GRP 1:v��Fr	v���+�+��߇�?(OCDO[[ ���@hp�fhp^EZOlL �� ߢ�6�?�O�O�OPOrOX�O�E�!MR�3�=T֏���ra_s^�_�_�X_�_|_���!OAD?BANFWD�/�#{ST�11 12%�`  4OSSW)���ߣ�B��B�p�L��D��3EɚƑ5^hFrto�F\o no�o�o�o�o�o�o�o �oC"4yXj���������r���mmh�o�p��[���ex<�N�
X0�B� T�f�x���������ҏ ����M�,�>���b� t���������Ο���J	g2l�$b� ߯ �[������֯��ǯ ����B�!�3�x�W� i���������ÿտ� ��"��?���cϨ� �ϙ��Ͻ������� J�)�;߀�_�q߃ߕ� �߹���������*��c3C�U���<���H	g4r�����	g5��������	gA6�*�<�N�	g7k�}�����	g8���������	gMA�P��N�  	dOVL/D  F��O��	dPARNUM � k���hS[CHc	 q�p��#UPD���d��_CMPa_�0-�3 0' e~|ER_CHK��� aB����RS?P�_�!_MO��_�_���_RES_G` F�E`Y/ M	e/j/�/�/�/�/�/ �/�/??=?0?a?T? f?�?�?�?�?�?�?O �?O9O,O]OPO�OtO �O�OK=#B�F/�O�O __>_1_b_U_g_�_ �_�_�_�_�_�_o	o :o-o^oQo�ouo�o�o �o�o�o �o$)LZ�O_Gq��L�O g;%�����=#� ���=#j��!�&� =#��A�`�e�=# ��x����="V 1!��+�  �[�J؄Y��T?HR_INR$ h��d�d�MASmS$� Z8�MN#��V�MON_QUEUE "��+��8��N�U�N8f�����END��%/�řEXEԟŕFB�EӐ���OPTI�O��.+��PROG�RAM %��%���ޏ���TAS�K_Ie�OCFG #���}����DATA_ 1$���@+>+� 2 ��� ���=�O�a�k��  ��������p����ѿ� �����4� �������  9N����h�_��q�{�ܯ�ϭ��9 @Ұ��������߳�g�/�A�M�^�p�㬏INFO��X�2� ��]���������� � 2�D�V�h�z���� ��������
��.��ׂ��&���Tx��K�_��'����p�ECNB(�8!��2��ں�G��2(� �X,		�=������@�  $� �		� ���6l*<�p��_EDIT )�����WERF�L���#RCRE�P *�� B����9 
�̯`�
M�P�RGADJ +�
A<�?�4����z�,����?�  BzD��<v��%|`/BT|���2.�V�	H�@lE{�Bh�N8�@\��-*� /�" **:�"�/�&�/�Gy$P�8� �/� /?%8�	���/?a?o?-??>Q8gr_?�?�?�?�?�?�?9OGOO2?>y$ЀA��/_O@�OkO}K��A�AЀ {M�O�O�OU_�OQ_;_ 5_G_�_k_�_�_�_�_ -o�_)oooo�oCo �ooyo�o�o�o �o�oqmWQc ������I�� E�/�)�;���_����� ����!�ˏ���� ��7���s�m������ ��ߟٟ�e��a�K�E�W��H	O��<���t$ 3�E� �h������l#x$�'�����C� �/�/�/ů{�ͯ���� ρ�+�}�g�a�s��� ����������Y��U� ?�9�K���o��߫ߥ� ��1���-���#�� G���}��	���� ������u��q�[�U� g�������������M ��I3-?�c� ���%�! �;�wq�� �����i//e/ O/I/[/�//�/�/�/ �/A?�/=?'?!?3?�? W?�?�?�?�?կ.Oq� >OdO/��OS��OGO�O��O�3�$PRGN�S_PREF }/E�԰�԰
ñ�AIOR�ITY  �4��R��AMP�DSPON  d��İ�EESUT-V���Q+�AODUCT_ID E�8R�O�FOGGRP_TGL-T�V�V�HIBIT_DO�LX�[TOENT �10�Z�@(!AF_INEkPo)g?!tcp)oQm�!ud@oyn!icmho�m"R�OXY_CFG �1k �ӱ)�� ���o�o԰� �o�eD+hO a����������@�R�*�S�b	3
Y[R% O����B�?���6��/̄����4�SU���A���,  �P�Q�c�u�OX�f�Z鏸�ʟܟ���3g�ENHAN�CE 4s�#�A≛d�N�5�  	ʰVT5
_T�a�A�PORT_NUM�-S԰8U�A_CARTREPLP|�l!RSKSTAkW��[SLGS`6�k�1�ӱUn?othingV�7� I�[�k���������_���TEMP 7�Yÿ�5�_a_?seiban�O&� �O6�\�Gπ�kϤϏ� �ϳ�������"��F� 1�j�Uߎ�yߞ��߯� �������0��T�?� Q��u�������� ���,��P�;�t�_� �������������� :%^In� ���� �$ſ>��VERSIJP�W�_ dis�ableh�;SA�VE 8�Z	�2670H7955!�!>���zo� 	(uR�?I+	@/8#e]/�/�/�/�/�*u,��/��z]_�P 19k� �\m�D2�L��7V?h?��^�@URGE�B�P�^"QWF�0�Q/T#���VW`�4����WR�UP_DELAY� :ʭ�eWR_?HOT %~�wR�=�-O�5R_NORMALH8ROqO@GSEMIPOvO�O�A�QSKIP,22;~�=3x�O_0_�B_]~�i_wWQ�xs�HP_�[ 	#���
C�_�[u_�_ a_o!o3o�_WoEogo �o�o�owo�o�o�o �o-SAw�� a��������=�+�a�s������$�RACFG <��K!�8#���_PoARAM�A3=�Kw @ �@`�6�#�2C.��1"&��C�6��B�����)�q0��BTIF���:��CVTMO�U�ѥ���D�CR,3?�IE0��QC˔�E�i�EMU�D���2!B�L�]�P���a�8%���tA�{qE�_%�Q_ ;�~��;DAP���g;�-�<�A7���!������P ��¯ԯ���
��.� @�R�d�v�������� п������*�m�N� `ϣ��ϖϨϺ����� ����&�8�J�\ߓ��DIO_TYPE�  3=K�a�ED�PROT_��@��Gʐ8$B�SE�*����BA�� �H�B�6���H�:� �^�I��m���O ��Y_��M����U� C�y�g����������U ������	?-O Qc�������{ �;)_M� ���{�w/� %//5/[/I//��/ ��/a/�/�/�/!?? E?3?i?�/�?�?a?�? ]?�?�?�?�?OAO/O eO�?�O�?mO�O�O�O �O_�O+__;_qO�O��_�S��INT 2�BEVE��рy�G;� �_�[%�E� or�f�0 o0kM_Po A_`oboto�o�o�o�o �o�o(L2D �p����� � �$��H�Z�@�~�l� ����Ə؏����� � �0�V�<�z�h��������FPOS1 2�C~�   xAtHome	o������Q��a���f�uſ��ؾ���m�<���5/��5?� � G���AtPOounc������d�o3�A�S�Y�R	3����{������ï4
����|��$)�;�5����k��� ����K���AfD��� �!�3�E�W���{�� ��������^����� ��A߬�e�{߉ߛ߭� ��H���i��R�+�=� ��a�s�������� ������'���K����G�
AtMainOtPsn���� ���,������TipDOress2��Ф?QK���nu�als Chang`�������K�AtAuto��ٶ�/AK�&Y�urnֹ�/(��K�q2/�����//1/��	[*����s/�/�/�/K�aj[.����/t?? !?K��[/ڵ�c?�?��?�?K���Pos1�?ٶ��?dO�?O#OZ/׸�SO�OwO�O�O	sկط��OT_�O__sM�ط�C_�_g_$y_�_sſط��_Do��_�_os6Joٶ�`3o�oWoio{os7�o�ٶ��o4�o�o�os	8:ٶ�#�GY&ks9�ٶ���@(��L��u�4@0U�ڵ�;���7���͉2 2DΟ���� 2���9T�u�{���� :�\�ҟp�������� >�ܟ'� ����6��� Z��~�鯢�į:�د ����� ���D���h� z�Ϟ�$�¿K��Q� 
�,Ϣ�@�R�d��ψ� ߬�������k�ߌ� *߳�N߹�rߔ�
�� ����U���v��_�8� J���n�������!� ����r��"�4���X� ��|�������;��\ ����Bd�x ��%�F�/ �>�b��� ��B/��/�/(/ �/L/�/p/�/?�/,? �/S?�/Y??4?�?H? Z?l?�?�?O�?�?�? �?sOO�O2O�OVO�O zO�O_�O�O�O]_�O ~__g_@_R_�_v_�_ �_#o�_)o�_ozoo *o<o�o`o�o�o�o�o ��C.g]�Y���ԏS3 2�E독��oO�:�<��5i�{��'�9� ]�㏁�̏����@� ۏa�����#���G�i� ߟ}�����*�şK�� 4�����C�ɯg�� ������ѯG����	� ��-���Q���u���� ��1�ϿX��^��9� ��M�_�q��ϕ�߹� �����x�ߙ�7��� [���ߡ������� b��߃�!�l�E�W��� {����(���.���	� ��/�A���e����� ������H��i� +�Oq���� 2�S�<'� K�o����� O/��/�/5/�/Y/ �/}/�/?�/9?�/`? �/f??A?�?U?g?y? O�?#O�?O�?�?�O O�O?O�OcO�O�O�O _�O�O�Oj__�_)_ t_M___�_�_	o�_0o �To�_do�o%o7oqo��omo�o��s4 2F��o�o�_l�_� o�O�s��� 2��V��w��Q�9� K�ԏo��������� ۏ�s����5���Y� ߟ}�������<�ן]� ������C�U�ۯy� ���&���G��!�	� ���?�ſc�쿇�� ����C��j�ώ�)� ��Mω�qσ�ߧ�-� ��T���O��%߫�I� ��m��ߑ������� ��t���3��W�� {�����:���^��� ��Y�A�S���w��� ��$������{ �=�a���� �D�e�'� K]��
/�./� O/�)//#/�/G/�/ k/�/�/�/�/�/K?�/ r??�?1?�?U?�?y? �?O�?5O�?\O�?WO O-O�OQO�OuO�O�O _�O�O�O�o|_g_�_ �o�___�_�_�_oz5 2G%�_�_�O �o_�o;_�olo�o�o �o(�oO�os� 2nVh���� 9��4��
���.��� R�ۏv�����֏��Џ Y��z����<���`� r��������C�ޟd� �>�&�8���\�⯀� 	����ȯگ`����� "���F�̿j������� )�ĿJ��q��l�0� B���f��ϊ�߮�4� �����ߑ�,߲�P� ��t��ߘߪ�0���W� ��{���:�v�^�p� ������A���<� � ���6���Z���~� ��������a���  �D�hz �' �K�l
F.@ �d��/�/� �h//�/*/�/N/�/ r/�/�/�/1?�/R?�/ y??t?8?J?�?n?�? �?O�?<O�?O�?o �O�O�O�_�O|O_�Ox_;_1j6 2HBo �O�OO�_4O�_XO�_ �_�_�_�_Eo�_loo �o+o�oOo�oso�o �o/�oV�oQ' �K�o���� ���v����5��� Y���}������<�׏ `������[�C�U�ޟ y�����&���!���� }����?�ȯc�鯇� ï����F��g���� )���M�_�心�ϧ� 0�˿Q��+��%Ϯ� I���m��ϑ��ϵ��� M���t�ߘ�3߹�W� ��{ߍ���7���^� ��Y��/��S���w�  ���!���������~� ���=���a������� ��D��h�' cK]���. �)���#�G �k�����N/ �o//�/1/�/U/g/ �/�/?�/8?�/Y?�/ 3??(_�?�?�?�O�?��?"O�?OXONZ7 2I__�?O-?�OQ? �Ou?_�O_�O�Ob_  _�_$_�_H_�_l_�_ �_�_+o�_Lo�_soo no2oDo�oho�o�o �o6�o�o
�. �R�v���2� �Y��}����<�x� `�r��������C�ޏ >�����8���\�� �������ȟڟc��� ��"���F���j�|�� ��)�įM��n��H� 0�B�˿f�쿊�Ϯ� �ҿ�j�ϑ�,ϵ� P���tϰϘϪ�3��� T���{��v�:�L��� p��ߔ���>����  ���6��Z���~� ����:���a����  ���D���h�z��� $��K��F
� @�d���� ��k�*�N �r�
/�1/�U/ �v//P/8/EO�/�/ �/�??�/??�/<?u?kJ8 2J|O?(? J/�?n/O�/(O�?#O �?�?OO�OAO�OeO �O�O�O�O�OH_�Oi_ _�_+_�_O_a_�_�_ o�_2o�_So�_-oo 'o�oKo�ooo�o�o�o �o�oO�ov�5 �Y�}���9� �`��[��1���U� ޏy����#������ �������?�ȟc�ß �������F��j�� ��)�e�M�_�诃�	� ��0�˯+�����%� ��I�ҿm�󿑿Ϳ�� ǿP��q�Ϙ�3ϓ� W�i��ύ�߱�:��� [���5��/߸�S��� w� ���߿���W��� ~���=���a��� �� ���A���h��c� '�9���]�����
�� +�������#� G�k���'� N�r�1mU b?��/
?8/�\/��Y/�/�:MASKW 2K�;�"�/��'�'XNO  ¹/ �0?6�1MO�TE  �,�4/1_�CFG L6=�c4�:PL_RAN�G21.!�5�s6OW_ER M�%�0��6SM_DRYP�RG %�)�%�3/�?�5TART �N�>�:UME_�PRO�?�?MO�$_�EXEC_ENB  w$�2f1� �GSPD&@h@pH=�7GTDB�O�J�RM�O�HIA_O�PTION�4c1��3�ANGVE[RS�A�*<O��)I_AIRPUR�0 .J�$c_�+MT_� T�04;�5�OBOT_ISOLC�,�_P`Qj=�R/NAME\�$_�\?_CATEG�(�3��#j2k3ok
cOR�D_NUM ?��8\QH799�j`869p`w$�zo�o�$PC_TI�MEOUT�? xު S232O21O��%�C LT�EACH PEN�DAN�`[f5f0��\2/0 KC�L/C @nce �Cons-"{�# No Use^}`r������"�bNPO� @�bf1�E�aC7H_L)@P�^d�	=��!UD�1:c�
�R� VA3ILSa�E�5Q�SMFST_CT�RL 3R�+D%���/ ߏ�"��^_E�4�i� l�1��������ɟ ۟���	�/a�4�� X�K�|�k���o�	�ϯ ����)�;��K� x�G���������俳� M��%�7�I�[�m�� U����ϋ���ӿ��� (�����W�i�{ߍߟ� ���ߙ��� ���$�� H�7�l�;��ߛ��� ����������D�� h�[��{������� ��'9K!�[� �W��������� ]#5GYk}� e�����// 8/�g/y/�/�/�/ �/�/��?�4?'/ X?G?|?K/�/�?�?�? �?�?OO�/'?TO#? xOk?�O�O�O�?)O�O __%_7_I_[_1OkO �_gO�_�O�_�_o�O m_3oEoWoio{o�o�o u_�_�o�_ �_$ Ho�ow���� ���o�o ��oD�7 h�W���[���͏ߏ ���'��7�d�3� ��{�����П��9��� �#�5�G�Y�k�A�{� ��w�̯���߯�� }�C�U�g�y������� ����쿻���4�#� X�'����ϙϫϽ��� ����ɿ�0���T�G� x�gߜ�k�������� ��%�7��G�t�C� ��߼�����I�� !�3�E�W�i�{�Q�� �������� ��$�� ��Sew���� ������� D3 h7������ �/�@/d/W �/w/�/{/�/�/�/ ?#?5?G?/W/�?S/ �?�/�?�?�?�/Y?O 1OCOUOgOyO�Oa?�? �O�?�O�?_�O4_O �Oc_u_�_�_�_�_�_ �O�Oo�O0o#_ToCo xoG_�_�o�o�o�o�o �_#oPotgo ����o%��� !�3�E�W�-g��c ���܏ˏ ��i�/� A�S�e�w�����q��� ؟����� ��D�� ��s���������ͯ߯ �����@�3�d�S� ��W�񯷿ɿۿ��� �#���3�`�/���w� �ϗ��ϛ�5����� 1�C�U�g�=�wϤ�s� �߻��������y�?�Q�c�u�������$RSMFST_�SV T��}����	����ӎ����}�	�&T)�H%�!�������MASH_ENB�  �� ��PR�G_ALRM  ���
�����D'SBL��)�����U��2�F�/	��/
��h/o	/��k��f���_CHEC�K V�MN�CON9���DIALM 3W��/�A=�"4�R�UN��M��SHARED 3X�� �����8��xTRBa��PACE1 3Y~�� 
�:C	/��j ��{,7<��?���/ ��/�/�/�/?	76/ H/Z/l/?�/�/�?�? �?�?�?�=����M:? L?^?p?�?�?�?�O�O �O�O_�O_2?HOZO lO~O0_�O�O�__�_ �_o�_2_D_V_h_z_ ,o�_�_�o�o�o�o �o"@oRodovo�o�o �o�o���	��� <N`r�6��� ��Ꮰ�����,�J� \�n���2�������ڏ �������F�X�j� |���@���ԟʯ믚� �!��6�T�f�x��� <����ƿ)��������2���!2",��4/ j�|���@ϲ����-� ���>��S�P��ϕ� �Ϲ�k�������O��� �L�3�a�ߑߣߵ� g����������'�H� /�]�{������u� ��	���Y�#DV= w���������q�� ��1R9g� ������	/ �-/N/`/7/��� ��{/�/?&?�/ G/\?C?q?�/�/�/�/ w?�/�/O?�?7OXO /OAO�?�?�?�?�?�O �?O_0_�OQOf_M_ {_�O�O�O�O�_�O%_ on_�_Aobo9owoT�3g�yϯ_�_�_�o �_)o,rob�Z��o4�o�o�o�o�o �JM��-�����{����5���� �Ǐ9�k�n���N���ş��ڟۏ6� �� $�6��Z�����՟o� ů毽�����7�!� 3�E�W�	�{�������@����޿��80� B�T�f�x�*Ϝ�ο�πϱ��(���=�>�Gw ]T� 8�:R�
�� �߷� V�T���������,� X���I�x�V�u�ߨ���d���������� �+�=�O�E�W�i�Z� ������������S� /ASe[�m���� ������
��s= Oas�{������ `9� @��%��,/_/( /��/�&�!�x# �/�/�/?�%�/ ?B? T?r?(?Z?�?�?x?�? �?�?O�?�?�? ObO tO�OHOzO�O�O�O��
L/_�k_MOD�E  Tɔ�6VS ^T�_��A��H/q_�_�Z	�_�o�dCWORK_�ADC\�(�^�aR  T�a��Z`oD`_INTV�ALCP�Đ\�lfO�PTION{f ��e�pTCFq�_�T���İX��c�bV�_DATA_GR�P 2a�_�DP�_(�_L7y �Oyg����� ���	�?�-�c�Q� ��u��������Ϗ� �)��M�;�]�_�q� ����˟���ݟ�� #�I�7�m�[������ ��ůǯٯ���3�!� W�E�{�i�������տ ÿ�����-�/�A� w�eϛωϿϭ����� ����=ߢi�8 ��\B� ߮������ ��,��P�>�`�b�t� ������������� �L�:�p�^������� �������� 6$ ZHfl~��� ��� 02D zh������ �/
/@/./d/R/�/ v/�/�/�/�/�/?�/�*??6?<?N?�?���$SAF_DO_PULS.`�`	q�c��1�0CAN_TI�MBQ�S�f�1R� b"��"6�PP��P�P
�T	��R�Q	C�Q�1�R  ��3OEOWOiO{O�OO��O�O�O�O�O_W�(	q&P�R24Td �4�1?Q?Q;U�B]SY @�o�_v_�_�#R�1�_�WP�U�"'�� tP#RTY`0P��_o#o5o?fT D��?ohozo�o�o �o�o�o�o�o
. @Rdv��_�Uu_�����r � .R�P;�o� T��Qp�4�v
�?u��Dk@�A�A�z�� � �B�Q�QA�L�D�1 �1��������Ώ��� ��(�:�L�^�p��� ������ʟܟ� �� $�6�H�Z�l�~����� ��Ưد���� �2�D� S��_o������� ��ɿۿ���N��R#� /�A�S�e�wωϛϭ������#R0�RY��U �Q�1 UAw�k�6�H� Z�l�~ߐߢߴ����� ����� �2�D�V�h� z������������ 
��.�@�R�d�v��� ������������� *<N`r��� ��%���&8`J\n��Y��R���1P� ��R��}�� �����A� ����/#/5/G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?OQOcOuO��Nc�O�O�O�O�O __)_;_M___q_�_ �_�_�_�_�_�Z��_��_#o�t��t��o�}	1234�5678@�h!?B!��
��
/��@ �o�o�o �o�o�o�o!'q�O J\n����� ����"�4�F�X� j�{�9����ԏ� ��
��.�@�R�d�v����������}�BH ϟ��	��-�?�Q�c� u���������ϯ��x����:�j#� M�_�q���������˿ ݿ���%�7�I�[�mτ�D�wϟϱ��� ��������/�A�S� e�w߉ߛ߭߿߂��� ����+�=�O�a�s� ������������ ���9�K�]�o����� ������������# 5GYk*���� ����1C Ugy�����D�f���/-/l?/[jC�A��J_   ��H2�B� } ��L&
�'�  	�bb2��/�/�/��/	<�O
,��`1� 3 4bb  L2T?f?x?�?�?�?�? �?�?�?OO,O>OPO@bOtO�O�O�O95��B(bbP�D�O�O�O_  _2_D_V_h_z_�_�_ �_�_�_�_�_
oo.oD]hbb
!�!~"<\d� Re�!  �lk�o�Fib�!>�!t  s �i��o9h`Z!�$SC�R_GRP 1d�"Y�"b�� �� �Z!� y%	 /q�r*r #t!Kc:wK6wdR��O-�� �rD��p��=0s�w�{�-<M-900�iB/700-IF 67890� ��t[qM9B7���C
V09.�00 9�Yx1q�+ ]�q�Fq hsq-3[a�q'z\qn�	_���ɏۏ���~���H�p���wx� H���D�1�Đb�6C%M|=��o� �(.�R5q�X���4��'
�"���²�O���5!�  ==��D�2�M�LCG%W(p�/Z!��̟��Bh��CY#hz\ ,UyB�  9��K�5qAs a�  @[ y�]���?e ��5��a ����5qF@ F�`ܢ�۟�� ,��<�b�M���q��� -�y���տ��ҿ���B�ϙ�J�5�n�Y� ��}Ϗ��ϳ������ ��4�F�,>�stf׋߂y'� �߽�Y"��@�e =@�w%��6p@�p��K���12345�#���$S�DA�wq�"��*Zsf`,2K�Z! ��C��g������� p�	�����E @��OW�i�,ߍ�x���.���x /��<��s��r/p ����p�f&r��8y?8��cN?W�8������R��sSV�GUN syst�em 0�	� �)�-�[vd]�N so�r�-3����塏�������/7�H���(�;�@/S{�G�VL/v/�/��/ ���/T�/�/�?6� @?Z�y�e?����?�� ���?�/�??O�?*O ONO9OKO�OoO�O� ���O�O�O�&_�OJ_ 5_n_Y_�_}_�_�_�_ �_�_o�_4oKߡ;/ ��ߨr�߷o�o�o*9 ��-� B�Of� �/p������ ����=�O�a�$o��p�����d��/���$SECLV�L  ���<��j7��L_D?EFAULT�����HOTSTR%��9��MIPOWERF���1�_�WFD�O&� 1� ��RVENT 1e���R� L!D�UM_EIJ�̙��j!AF_IN�E%��`t!FT$�����=�!tZ��`v�,���!RPC_MAIN���l��x�կ��VIS䥯k��į!�!O�PCUA"�H���m�!TP`�P�Ud�әd\���!
�PMON_PROXY��֖e��π��ӿϝf��Q�!R�DM_SRd/Қg@ϝ�!R5��ԘYh����!
��M��Мi��5�!RL�SYNC6�\�8|$߁�!ROS�����4p���!
C}E��MTCOM�߲֖k���!	��C'ONS�՗l�e��!��WASRCdl�֖mT��!��'USB��Ԙn����!STM���Қo��I�P�m�`�:������ICE_KL �?%�� (%SVCPRG1��D����2������3D��4.3��5VD[��6~���7� ���&���9������#����K�� ��s�� ���H� ��p���/��� ;/���c/���/�� 9�/��a�/��? ��+?���S?��/ {?��)/�?��Q/�?�� y/�?��/O�/�� �������fO�O�!�O �O�O�O�O__?_*_ c_u_`_�_�_�_�_�_ �_o�_o;o&o_oJo �ono�o�o�o�o�o �o%I4mX �������� 3�E�0�i�T���x��� ��Տ������/���_DEV ��?�MC::�L�?GRP 2i��t����bx 	�� 
 ,��t�. 7�����ϟ�ȟ�� )�;�"�_�F���j�|� ����ݯį����7����k�D��t��� ���������ۿ��� <�N�5�r�Yϖ�}ϏϠ�ϳ���G���t�  ���0�V�=�z�aߞ� �ߗ��߻���
���.� �R�9�K��o���
��(t������� ��6��Z�l�S���w� �������������D+h�a� x�	X����� CU<y`� �������-/P�-�b//�/m/�/ �/�/�/�/?�/?:? !?^?E?�?�?{?�?�? �?�?��OO�?AO(O eOwO^O�O�O�O�O�O �O�O_ _=_O_6_s_ Z_�_�_ O�_�_�_o �_'ooKo]oDo�oho �o�o�o�o�o�o�o�o 5Y�_N�F� ������1�C� *�g�N���������������ޏ�qud ��R�"�6 2� 	�T�3�B�����bO�A��1�����'��qY� ����A��r�-��:b���:y��B�\\�?����@�;A���@H�+A����X�%JOGG�INGX���R��=�i��{z�?����-��>O~�@��d���U�����1�i��6Β?D��vAq�����(?�0@5��1��O�����)�����@�����m��V��1�>�2x�����AV���@�6�-(?�u�1��Ư��(�6�i��9�z�8b�?2�;�N40���G=����1�����Mi�@�">�G�5��U�K�hY�g��!A�a���7@�;��u��b�M]1�?�S�5@��?�� �@��Q�eZ˿��F��ػ���ߡ)��?���������(�D콈�/���̿u�1����T@AZ}A�1�KjA�p@&�Y��~>ʌ����@nn�i�!�" �1��@=@�@�Pj�A�K�AW�����?���}���tϳ�<��@;������?���>��������X�����WA�AI�.���~Aw����r�Y�f�� �C�u�%�,A�yP���)��F@��9�����?�A!��?՚A�}�Q�c��H߳�깶�1����?N�=��%�$`B���}1�����A$��A7?����aA�u�)�;�1�A`c��%7nA�p*���>� �)�O�L@�������@v�w����oA���%�7��ߡ�1��u������?����2��R����81�=(���A��Ap��� P�An�@=�քY��f<�l���@\�9��u^­���4��kU�;7�@���h�C[�A��x��'7���C������/⩹��C�;���>��l=k�U�r���1���"�g]qA,z����rSAch��@#x�Y�w���̉������j����^nU�����@���r)�@���]����?�z�����,��奿��� ��?!��2�!��ؿ�n>�lPU�����AW��A5�}�h�AY�N��Q���G��!���=���j��|��!��W��?�S^����A5������Z��������ߡ���w-���	?r"->��mƿn����F���w�A�q�\A!��� �Ac�x@�ec5Y��}�����Q���D���I�����v,�)�f�J���ϑLi�9*?�уu�l��	���^j�~�>ʜ�>%��[��S?��پ�\	An���AJ���&I�PK_������VM��a����+���u�i)�*�!�@FEY�|VH�AN�#���?�y�I[@/��t�2��@B�;�g^�C)��B���� 7�@�=�A��{�����Agn��}������}E�@�1���g���A�q���n��$�B?^/-/?�����`�^�9���k�?��@N�`��6������,��/��Aj8�@M�e�@� H@�����.FA�x����������±-T�ZL�)�Gm{��AE����@����ٿ/ ?�?���Y)�<N9��D�a"�.�� �f^1�`�>@/�ƠAXl����D3Ad�����dY��(���;��?�:+��w��1���^ǁ��!��A�P�Axn���k�A��$�?8�?�O��n��A�����9�h��q/���2�A�����a�A6�^��}��'߿�ݧ�g�:V=�������]�U����PA�@����A9^h��?�Ab�`�O�Oܐ_��Sa�@����w�?y�N�I�A�=�c�پ�@ΉcA����c@���}@F�sY���mi�3�U�l���9lG�¬��J��JT��!��7U@r�A��Ib��2ᾨ��<m__do����;�|}�,e��@8�I��OV��	��پ>A���@�̈�4��@4+�@8���Y���^�j�����ӟ87a��¤���e"��)���@��?@�8�Aō�0@*�@U��AjTD_PO�UNCgo:|y`]���l���=m�@ �iI���"��z�پ���_A&S�@>@� �?��@Z�J�Y��J�qh��(>9zb���E@� ���o�`��S@���gA��@����?mG"�Fv��B�� "@U��¿	�V�\�h�>�W?����U��R��^�#A,
h��wt�QIӡ.�	ӨA�u����?�;<����1�BQ4����Ed��ZPA����A1aAg����o������G��:��?��-a�`wВ>'�ʧ>�u��@!����iW�A>�GQ�L�'��T�Wm��kA������P;?��#:xBP����5��V�h�A�wA\?��A�Ƌ��ˏ\��Gt���2�"������d?�'9���n�>	q/)Δ���?�P�@����G�qBI5^�� &С.C��A�ͅ�6=D�;�@�1��BY.�)��w�@��Á@���@�A�¿��sBvܑ�CC?_AUT01����ߗR��\���j����'??�>I��G�7���:��0@�	��A0������@�@%:�t
9�����c����D�:��D�haJ�����)�z�@�w�@�&�8A� ��%@2]"AoSo\��w`����E;,}RA��V':�@��ާ��`?g�qNR�ZAB;|�AICm��SAfD3��{h��3��������v>/���m+���A��߿׵�6A��3`�2���2&Aß�9�K�0�o���E��@ua��g�b::��\� ���)�qN�g�f��A�PK�0o�_A�r��]�M��4���-���c>0�/�l;cᰩM>:���j<�=�A������mA�~���o�ݥu��
�Y�;R�V'��D@�T�)����@A?AR{�EAA������4���'���� >0S������|\�M>�[�A0^o���N%A ;��Pi�I`��������o��I�|gbN1��U�z�VG��r!����A4�V��V!e��4M��������b>0fz±߿%�}0��"��P@׏��1�
�A%M������}�ߧ�j���QvZjW�a���?�Q=�V�x`��Y�J�Y2}AX��A˞@x�A+�(?�8��]�)$����l�����>O��°U���L�|�2`@����2��s���k�A@`d�����o���*�x��_�vG>��<���߾�J����uM��@���@^[C��|O���@h��.9�����1�6�#;�=� ��¯;�BP*���"���AC[��AnfGA��H?�}n]�o�T���8�E>�wg���0�>eI<�9����Bܾ�T~%M>�3@���	@j�+������2�@u5�������E��'��=ș��¯3HBPW���(�,@��W�A?I�Ad]��A���?Gu�1C(��f�Io%���p���Q���\�zqN(��@�«�A�@o�п�p?�?���C>�M Q�<sH�A����¦�rA�ӊ�!N��?�Ӽ�A:���J�d�A@��@��y����rY)�(����A]�;�:&�����?�@�
�A� �Q�����@���>���M!@<f�߱A�����A���qnr�h�`�A�\c��M��A3 ?�@�p���/w`�^|͐�I�<��@[�ߪ?����R�
�2>y���1����^�AFh{3�N![���6@���wB-A�4�������J����¬#���=@�������c��ua����4�	S012�SSWy��=,R����%@�0s?�!�;>���;�w��}.�>�/?�ҧ�
���@�� �WSQ�@��ͨe��pQD��PC��2�پ���³�~��/������T�@z���+ɇ��o�̎?sOsc^�S�Qv#P�?"س�%:��1ѿ�$�����=�o�`'�qAo�"�n�AO�ja�Q,^�������@��7!ua����[f-O?@x���A4k5a����Ai���*
_�ALTMASTE�RzONZ$S ���%<%#��8�]�Oer�5���Y(Z�
��N��c@���A���=� �A�ݴ��;t�;�D��,��B�X_ ^?�p@�p�#AC��@���?A���@�r�jq�o$�S�Qv�v>�J�E@Y컳�F��%O�!����� P�A$ʿ6@�����Y��L@.?�`����k$���z���£ٌ��gj��{�@���h@�W�A����@?��@���RETHOM�"o�l5`.���[�%!�.�]��Z���"��9q�A��AF�s�=-��?�"༪_�ª��l%���"��2�£�g�l���e���]S^�?
`�A�~�@1�)}�/�%5`3%���\:�!!�yE����LA �AE��u�>�?��`�=r�oZ��l'��W�{upvyp����" ��L@����A���
�^�u/����r�Oc�%��S?�S�¿n;���>�\�?�'��Q���a��z�KA���"?��1>N A��EhA�\���%H.9}��B�nB���Q��W��*��A����@���A~���������p� SP0�A���<?l"߸��{35�>�ߋx?Fz�?���I�]zEA/���K�h�@����­^	��BA�/z����n��d��FXB]�XY?@���8�P7AQA�A�'ı�_MOV_�`Er��F�	��Em�)���!����,�9��>���-�(���0���A7����S�Q�N��@1����^
PA�����������7B_?}��Ivp@3���7�Ah0OA�Ƌ@�������POA���+x�& %��{A�^��Ơ�G�A�#:���~`?���џ��A�݅�������5�B_9`��� 4@��l�@���Af�e�A��ſ�y������+�k1����=�b>
����@;�Ia=�O���^�����o� @�>L��PK_���0���y��A�?����ڽ��Z�H�B]���%�W��Kd�AR��@��M��!�3���W���A����=*�� ��<N5�<�an=	q������f��A9����~�5�U��,B\�ݓ��A���`��P�����V;B�]0}ՎF���Q��A#ެ?An~��,Z���~�ȉ�l��^Ļ��v���X�����6�A/V!��:���*����:�!ߺ�A��-��R)���YA��FE�}����@����A���A�1��A���@�v�~�c�~����LS�8=�μ���;���=@��?����^���A3���~���:R��/�A�A�gi�������wf�oB\�aI�F9�����A
��A�x9��S�8��2 �y}ye�S���w���������%�>����� ?-cQ�u��� ���;) _M����s� �/�/7/%/[/� �/�K/�/�/�/�/�/ �/?3?u/Z?�/#?�? {?�?�?�?�?�?;? O 2O�?O�?SO�OwO�O �O�OO�O7O�O+__ ;_=_O_�_s_�_�O�_ _�_o�_'oo7o9o Ko�o�_�o�_qo�o�o �o�o#3�o�o� �oY������ �aF���y���� ����ӏ����9��]� �Q�?�u�c������� ϟ���5���)��M� ;�q�_������ί� ����%��I�7�m� ������]��Y�ǿ�� �!��Eχ�lϫ�5� �ύϯϱ�������� _�D߃��w�eߛ߉� �߭߿���7��[��� O�=�s�a������ #���3���'��K�9� o�]����������� ���#G5k�� ���[����� C�j�3� ������/] B/�/u/c/�/�/�/ �/�/#/??�/�/�/ ;?q?_?�?�?�?�/�? ?�?OO#O%O7OmO [O�O�?�O�?�O�O�O _�O_!_3_i_�O�_ �OY_�_�_�_�_o�_ oq_�_ho�_Ao�o�o �o�o�o�oIo.mo �oa�oq���� �!�E�9�'�]� K�m��������ޏ� �����5�#�Y�G�i� ��я������ן� ��1��U���|���E� g�A����ӯ	���-� o�T������u����� ���Ͽ�G�,�k��� _�Mσ�qϓϕϧ��� ��C���7�%�[�I� �mߏ������ߵ� ���3�!�W�E�{�� ����k���g������ /��S���z���C��� ����������+m� R���s��� ��E*i�] K�o���� /���#/Y/G/}/ k/�/��//�/�/�/ ???U?C?y?�/�? �/i?�?�?�?�?O	O OQO�?xO�?AO�O�O �O�O�O�O_YOOP_ �O)_�_q_�_�_�_�_ �_1_oU_�_Io�_Yo omo�o�o�o	o�o-o �o!E3U{i ��o����� �A�/�Q�w����� g�я�������=� �d�v�-�O�)���͟ ���ߟ�W�<�{�� o�]������ɯ��� /��S�ݯG�5�k�Y� {�}���ſ��+�.��. 	� 
 U,�.�.�.��&�� �K�2�� sυ�lϩϐ�����B� �����5���8�b� �φ�mߪߑ������ �����1�C�*�g�N� ��r���������	� ��?�&�c�u��ߙ� P�����������) M4q�j�� ����%|� [fx��� ��/�3//W/i/ P/�/t/�/�/�/�/> ??�/A?(?e?w?^? �?�?�?�?�?�?�?O  O=OOO6OsOZO�O�O  ?�O�O�O_�O'__ K_]_D_�_h_�_�_�_ �_�_�_�_�_5ooYo �ONo�oFo�o�o�o�o �o�o1C*gN �������� �ro?�Q��u�\��� ����Ϗ���ڏ�)� �M�4�q���j����� ˟ݟ4����%�7�� [�B����x�����ٯ �ү���3��,�i��P�����d �R��!�{ 2 	? � ݣ��м���@���пӿ���M������9 �G�%�G�lϨ��R�"�6��?V�?����Ϝ�ǹ���p�ϧ����c����B������%TD_G�UNs�F�>R��,����cތ���@ֻ�y����K�ߣ���?�����JOGGIsNGF�t��É��:���������I�O�MS<q�w�Bу��� Z��﫰��Y���������B�#�C�V>E�K�CiAim���������������!����]�?����A���,����ź:�D���UU��1��JoTf���9�?������,��Ci� �E*/i��{ ���>��/����bvm/s/����ȕ/�/B���f�/���?)� ��]�t���/�/�2��.A?G?Š��<i?o?�7�6�?�/h�/�?!4�)7�V�?��?� �OO����=OCO�GH�}eO�?�?�O)�!G�]ֆz��OkO?����O�O��a2<__�Ns�9_�Oh�O�_�DJ)7wa_�?_�*���_�_���? �_�_�=?APog_y_^o�DW]����5oo@�;y�o�o��wZ�o�o�-z	�o;oMot2�Df]�O��	��o����ek��R7��Q_���}���;6������� o�c@�=�����/>f����݉��}/�POUNC�jތ�]!��,����@$7���yC�_:���ܨ���ȏ��섿B!�?� ���c��� y����VxM	��@��u1�����p�����@#�>�(��>6����쵯����V'ݯ�@��,��_�q�V���{^|]�?-�����A�������0�'����@�^��ٿ�	S012�SSW01Z�.�,�R��]�@N�y��߿���]Ϟc��n{�ϋ�@�í�������^S!�Vz?�ϳ�?�[?5�'P�S]Y�_����D��3�RETHO�M���SOc�ye��d����?��o���Ŵ�y�-�3���/�U���E����SP��!��;�Y�`s|�����Ŵ��o@�t�N���u����!���,�Α��_���|������<����W�i�N���!�=r9/$��K#��7�#��@k A�+="�y) �SAwe��� /�=/�/�)/O/ =/s/a/�/��/��/ �/�/??%?K?9?o? �/�?�/_?�?�?�?�? O�?!OGO�?nO�?7O �O�O�O�O�O�O_OO 4_F_�O_�Og_�_�_ �_�_�_'_oK_�_?o -oOoQoco�o�o�o�_ �o#o�o;)K M_��o��o�� ���7�%�G��� ���m�Ǐ���ُ� ��3�u�Z���#���� ��ß���՟�M�2� q���e�S���w����� ���%�
�I�ӯ=�+� a�O���s�������� !�����9�'�]�K� ��ÿ�Ϻ�qϓ�m��� ���5�#�Yߛπ߿� I߳ߡ���������� 1�s�X��!��y�� �������	�K�0�o� ��c�Q���u������� �7�G���;)_ M�q����� �7%[I ���o���� /3/!/W/�~/�G/ �/�/�/�/�/�/	?/? q/V?�/?�?w?�?�? �?�?�?7?O.O�?O �?OO�OsO�O�O�OO �O3O�O'__7_9_K_ �_o_�_�O�__�_�_ �_#oo3o5oGo}o�_ �o�_mo�o�o�o�o /�o�o|�oU� ������]B� ��u��������Ϗ ���5��Y��M�;� q�_�������˟�� 1���%��I�7�m�[� }����ʯ	������ !��E�3�i������� Y�{�U�ÿ����� Aσ�hϧ�1ϛωϫ� �Ͽ������[�@�� 	�s�aߗ߅ߧߩ߻� ��3��W���K�9�o� ]���������/� ��#��G�5�k�Y��� ��������{��� C1g�����W �����	? �f�/���� ���/Y>/}/ q/_/�/�/�/�/�// ??�/�/�/7?m?[? �??�?�/�??�?O �?O!O3OiOWO�O�? �O�?}O�O�O_�O_ _/_e_�O�_�OU_�_ �_�_�_o�_om_�_ do�_=o�o�o�o�o�o �oEo*io�o]�o m������ A�5�#�Y�G�i��� }����ڏ������ 1��U�C�e���͏�� �{��ӟ	���-�� Q���x���A�c�=��� �ϯ��)�k�P��� ���q�������ݿ˿ �C�(�g��[�I�� mϏϑϣ���� �?� ��3�!�W�E�{�iߋ� �����߱����/� �S�A�w�ߞ���g� ��c������+��O� ��v���?��������� ����'i�N�� �o������ A&e�YG}k ������� �/U/C/y/g/�/� �//�/�/�/?	?? Q???u?�/�?�/e?�? �?�?�?OOOMO�? tO�?=O�O�O�O�O�O �O�OUO{OL_�O%__ m_�_�_�_�_�_-_o Q_�_Eo�_Uo{oio�o �o�oo�o)o�o A/Qwe��o� �����=�+� M�s�����c�͏�� �ߏ��9�{�`�r� )�K�%���ɟ���۟ �S�8�w��k�Y�{� }���ů���+��O� ٯC�1�g�U�w�y��� ����'����	�?� -�c�Q�s�ɿ����� ��������;�)�_� �φ���O߹�K����� ����7�y�^�ݥ���$SERV_MAIL  �������х�OUT�PUT�����@��RV 2�j%�  �� (�-�k��������SA�VE���TOP1�0 2k�� d� { 2��6�s�y���6���'A���� ��������/A Sew����� ��+=Oa s������� //'/9/K/]/o/})�Q�YP<���FLT_CURGRP���}���'IDX�  }%�� ���!�/�$�'NUM��'��
�$DISF�U� ���-ER�R� ��/1��%=0T�I7��#�0�$ON  �/�?%��!�SCH 3l}%��V���! ���1�+OD4�$KO]O ��OlO�O�O�O�O�O �O�O#__G_2_D_}_ h_�_�_�_�Yp2�_�_ �?OOBo9Ofoxo�_ �o�o�o�o�o�o�o >)bM_�� ����_��oo 1o^�Uo��������� ȏ�ُ���6�!�Z� E�~�i�{�����؟ß ��	���)�;�M�z� q������ԯ���
� ��.��R�=�v�a��� ����п����߿�%� '�:�E�W�i��ύ��� ������� �&��J� 5�n�Yߒ�}߶ߡ߳� �������4�A�C�V� a�sυϲ������� ����B�-�f�Q��� u������������� ,P]�_r}�� ������;( 8^I�m��� ����$//H/3/ l/y{/�/����/ �? ?W/D?/?T?z? e?�?�?�?�?�?�?
O �?O@O+OdOOO�O�/ �O�O�/�/�/_�/*_ <_sO`_K_p_�_�_�_ �_�_�_o�_&oo#o \oGo�oko�o�O�o�o �O�O�O"_FX�o |g������ ��	�B�-�?�x�c� �������oϏ��o�o >�5b�t������� ��Ο���ݟ��:� %�^�I�[�������� ܯ����	��-�Z� Q�~���ǯ����Ŀ� տ���2��V�A�z� e�wϰϛ��Ͽ���� ��%�7�I�v�m��� �����߻������*� �N�9�r�]���� ��������!�#�6� A�S�eߒ��߶����� ������"F1j U�y����� �0=�?R]�o� �������/� />/)/b/M/�/q/�/ �/�/�/�/?�/(?? L?Y[?n?y���? ��? O7?$OO4OZO EO~OiO�O�O�O�O�O �O�O __D_/_h_u? w_�_�?�?�?�_�?
o oS_@o+oPovoao�o �o�o�o�o�o�o <'`K��_�� �_�_�_��_&�8�o \�G�l���}�����ڏ ŏ���"���X�C� |�g�������� ���B�T���x�c� ������ү������ �>�)�;�t�_����� ��ɟ˿޿����:� 1�^�pϧ���Ϥ��� ���������6�!�Z� E�Wߐ�{ߴߟ����������$SFLT�_WAILIM � �����  �!�T�,��REC_GR�P 3m����q�X� x �ߓ��߷�������������5� �Y��ZN_CFG nq��]����r�k�2o�q���,B   �A���D;� B}���  B4��?RB21���������!�GLOGM7ODEO� �Z�?OUT pq�9�� L�f��PXRQST  B	� �����THKCN�D 2q�� (o�������r� ��"4FX j������� �//0/f/T/j/x/ �/�/�/�/�/?�/? ?,?>?P?b?t?�?�? �?�?�?�?�?OO(O :OpO^OtO�O�O�O�O �O�O�O _6_$_:_H_�Z_l_��RPT1� rq��P^��  ��W�@���N@7
A\�G
G��q��p��q��Y�Q�Q�Q���Q�_s�[2�XJNo`oro�o�o�T3<o�o�o�o��nMPRL�E �sB	*MPST�A�PuF^y2�k|�o�3��W�T DATA �x�Z�d P�% �>�P�b���,����� ��t�Տ������/� A�S��w�����^��� џ������+�=� � a�s�����Z���ͯ߯ ����'�9���]�o� ��D�����ɿ����� �#��G�Y�k�.Ϗ� �ϳ��ψ�������� 1�C�U�g�*ߋߝ߯� r�������	���-�?� Q��u���\���� ������)�;���_� q�����X��������� %7��[m B������ !�EWi,�� �����/�// A/S/e/(/�/�/�/p/ �/�/�/?�/+?=?O? ?s?�?�?�?l?�?�? �?�?O'O9O�?]OoO �O�OVO�O�O�O�O�O _#_5_�OY_k_}_@_ �_�_�_�_�_�_oo �_CoUogoyo<o�o�o �o�o�o�o	�o-? Qc&���n� ����)�;�M�� q�������j�ˏݏ� ���%�7�I��m�� ��T���ǟٟ����� !�3���W�i�{�>��� ��ïկ������� A�S�e�w�:������� �������ܿ=�O� a�$υϗϩ�l����� �����'�9�K��o� �ߓߥ�h������߰� �#�5�G�
�k�}�� R����������� 1���U�g�y�<����� ��������	��? Qcu8���� ���;M_ "����|�� /�%/7/I//m// �/�/f/�/�/�/�/? !?3?E??i?{?�?P? �?�?�?�?�?OO/O �?SOeOwO�OLO�O�O �O�O�O__�O=_O_ a_s_6_�_�_�_~_�_ �_oo�_9oKo]o o �o�o�o�ozo�o�o�o��o#5GV{�$S�GWTSTAT �y���uq��pdu_�SPDUP  �t
thpHC_CFG zuw��r�x ���}�� d g ����p_2  |ts�@`x�pGRP �3{uy�pxx� 	 �pt	������Ï����uxp����� 3�ΏC�w�v����� ����U�g������&� ��ӟ�n�5�g���?� Q�c�쯇��"���ϯ �j����)�;�M�ֿ���Ͽϧ��sITF; 3�| ��� V��	��-�?���Y����}Ϗϡϳ�?�ELML�r|uu�u ������s�߫�%RSR�߭߿������ �@�+�d�O�a����������ߐ#���W�i���݁��qpr�����w@�B�!�܆݁��|��_�HK 1}m� ��t���M HZl����� ���% 2Dm�h_�OMM ~�m߭L�FTOV_�ENB�w�u��O�W_REG_UI��frIMIOFWkDL��A bv�IMWAIT�8	�u-#OUT�v̰���/!TIM�u;��a/VAL6/ #_UNIT��&��LCc�IO 3�
�C ���/?? 0?kT?f?x?�?�?�? �?�?�?�?OO,O>O PObOtO�O�O�O�Or ���O�O	__-_?_Q_ c_u_�_�_�_�_��$�SU 3��,\övpq
bwae�*o��4o����   couk_o�o�o�o�fB?��o�o1C�WL�ERR 3��,� ��ߋ��� ���	��-�?�Q� c�u���������Ϗ� ���)�;�M�_�q� ��������˟ݟ�� �%�7�I�[�m���� ����ǯٯ����!�p3�E��^�TRY�u��!MISg�3��, �R�Uk) ̿����Fa{q�����®a��Ϯ��I��4�m�_�_IRD_�MAP  �+����_�MB_HD�DN 3����#  �o����e�� ���2�)�;�h�_�q����c��ON_AL�IAS ?e�+( he&o������ Sj��P�b�t��1�� ����������(�:� L�^�	����������� u��� $��5Z l~�;���� �� 2DVh ������
/ /./�R/d/v/�/�/ E/�/�/�/�/?�/*? <?N?`?r??�?�?�? �?w?�?OO&O8O�? \OnO�O�O�OOO�O�O �O�O_�O4_F_X_j_ |_'_�_�_�_�_�_�_ oo0oBo�_foxo�o �o�oYo�o�o�o �o>Pbt�� ������(�:� L��p���������c� ܏� ��$�ϏH�Z� l�~�)�����Ɵ؟� ��� �2�D�V��z� ������¯m����
� �ǯ-�R�d�v���3� ����п������*� <�N�`�τϖϨϺ� ��w�����&���J� \�n߀ߒ�=߶���������ߩ��$SMO�N_DEFPRO�G &����(� &�*SYSTEM*��� $JO��RECALL �?}(� ( �}�ߔ��������� ���%�7�I�[�m�  �������������~� !3EWi��� �����z /ASe���� ���v//+/=/ O/a/��/�/�/�/�/ �/r/�/?'?9?K?]? o??�?�?�?�?�?�? �?O#O5OGOYOkO�? �O�O�O�O�O�O|O_ _1_C_U_g_�O�_�_ �_�_�_�_x_	oo-o ?oQoco�_�o�o�o�o �o�oto);M _�op����� ���%�7�I�[�m�  �������Ǐُ�~� �!�3�E�W�i����� ����ß՟�z��� /�A�S�e��������� ��ѯ�v���+�=� O�a�����������Ϳ ߿r���'�9�K�]� o�ϓϥϷ������� ���#�5�G�Y�k��� �ߡ߳�������|�� �1�C�U�g��ߋ�� ��������x�	��-� ?�Q�c���������� ����t�);M _��p����� ��%7I[m  ������~�/!/3/E/W/i/���$SNPX_AS�G 2������!� � 0�%/�/�?���&PARAM ���%�! ��	�+P����4� ���� OFT_KB_?CFG  ��%�#OPIN_SI�M  �+2�d?v?�?�3� POT�APCOUPL ;2��+ �05 �;� �1�%�9�1�?�?�OO)I�3EQ�3��,oO~$RVNO�RDY_DO  �5<5�BQST_P_DSBP>2|�Ow+SR ��)� � & S�012SSW01� 231 3 C7K 1�O�NC�TOP_ON_E�RR�O�"8QPTN� �%kP��CURRING_�PRMB_�BVCNT_GP 2��%:1�0x 	�O�_ ��_�_�_o�_4oo89do'e��iot.�VD�PRP 1��)	0)a�1ko�o�o �o�o2/ASe w������� ��+�=�O�a�s��� ������͏ߏ��� '�9�K�]��������� ��ɟ۟����#�J� G�Y�k�}�������ů ׯ����1�C�U� g�y�������ֿӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� �)�;�b�_�q߃ߕ� �߹��������(�%� 7�I�[�m����� ���������!�3�E� W�i�{����������� ����/ASz w������� @=Oas����bPRG_�0N�T16�kR�ENB�_�S}P�34K["�UPD 1��KT  
��"?/Q/ c/�/�/�/�/�/�/�/ �/??)?;?d?_?q? �?�?�?�?�?�?�?O O<O7OIO[O�OO�O �O�O�O�O�O__!_ 3_\_W_i_{_�_�_�_ �_�_�_�_o4o/oAo So|owo�o�o�o�o�o �o+TOa s������� �,�'�9�K�t�o��� ������ɏۏ���� #�L�G�Y�k�������೟ܟן韵_IN�FO 1�-%�  5�	 ��P�;�t�_�  ϼ3��z����Ʈ��5˿'�:��"6²��c��4"��C����B�� A�M�� D��1�ĐbKC%�O0=��������'�E�ټ�����D��I':�	::�^B���c��L���p�[�����G�Y����ʿ�������SYSDEBU)G�. � �d)>�SP_PASS��B?P�LOG ��*�7!  z ���?�װ ��	�  �� �UD1:\|�-�~�o_MPC�� ��(��	ߴ���2����?SAV �����"������SV�2�TEM_TIM�E 2���8 � 0  �� �e������j ����e��݌�MEM�BK  -%�����B�T���X�|�� @d� ��І���������,��K� "�@��#� 5�G�Y�c�q������������� ��� '9K]o���e�����! 3EWi{��������//��SIK��H -�@��xh/z/n��>*�B  ��7֘��/ ����� W/�/��ߩ � 8�	� �
?R?d? �p^��?N�@ ��?��b�?�?���&`�?���� �ODOVOhOzO
 �u��U�O�O��O �O�O_ _2_D_V_h_ z_�_�_�_�_�_�_�_�
oo.o"/T1SV�GUNSPDf� �'q��Q`2MO�DE_LIM ����ΦqaZ`za����LeASK_OP�TIONE�!�u��a_DI_�ENB�  ��q��aBC�2_GRP 3�@!�qð���@C�0�/q:L/KfBCC�FG �{�d֩�v�?п�� ��
�C�.�g�R��� v��������Џ	�� -��Q�<�N���r��� ��ϟ���ޟ�)��E�D��w����f� �����ί��J!�+� '���/�U�C�y�g��� ������ѿӿ��	� ?�-�c�Qχ�uϗϽ� ���������)��9� ;�M߃�i�T��ߩ��� ����i�����E�3� i�{��[������� ����	���S�A�w� e��������������� =+aOqs �������	' 9K�o]�� ����/�5/#/ Y/G/i/k/}/�/�/�/ �/�/�/??/?U?C? y?g?�?�?�?�?�?�? �?O	O?O�WOiO�O �O�O)O�O�O�O_�O )_;_M__q___�_�_ �_�_�_�_�_oo7o %o[oIoomo�o�o�o �o�o�o�o!13 E{i�UO��� ���/��?�e�S� ������{�я����� ��)�+�=�s�a��� ������ߟ͟��� 9�'�]�K���o����� ��ۯɯ����)�G� Y�k�鯏�}���ſ�� ����ۿ1��U�C� y�gωϋϝ������� ���	�?�-�O�u�c� �߇߽߫��������� �;�)�_��w��� ����I�������%�� I�[�m�;�������� ����������3!W E{i����� ��A/QS e���u���/ /+/�O/=/_/�/s/��/�&� �$TBC�SG_GRP 3���%� � ��! 
 ?�  �/?�/(? ?L?6?H?�?l?�?�< �/�?�?�?O�?3OO�WOAOSO�O�D�"�#�~�,dj5�A�?�!	 HD����O�HD�A p�4_V�J��+R��MP__�G>�
==sQ?3337_�_�[Z#@�O�XC��� A`�_�_�_�^0�_�_�_�^@-oumda �?�o�oyo�o�o�o�o0�o!>M{?�1S� ��gq	V3.0~c	m9b7�3	*�p�t�"�WvR�7�q�V�� �p�}�  �
��  �+�zB�@ I�;�b�q��/������ Ǐُ����!�3�E� W�i�{�������ß՟ �����/�A�S�e��w��������8{A�	�1234567�8�@ԯ��I��ͷ���b�t�}�V�!J2�#��-}������CFG �F�%�!)���(��]�˿ ��  �F�Tʜ T�z�eϞ� ���ϭ�����
���� @�+�d�O߈�s߬ߗ� ���������*��N� 9�r�]�o������ ����2 ��1��� d�O�t����������� ��*<��`K �o�����/�/ �5#YG}k �������/ ///1/C/y/g/�/�/ �/�/�/�/�/?	??? -?c?Q?�?�?{4:�? �?�?w?�?�?O3O!O WOEO{OiO�O�O�O�O �O�O�O__-_S_e_ w_1_C_�_�_�_�_�_ �_oo)oOo=osoao �o�o�o�o�o�o�o 9']K�o� ������#�5� �?M�_��?�����ŏ ���׏����C�U� g�%�7���������� ��	��՟?�-�O�Q� c����������ϯ� ��;�)�_�M���q� ��������˿��%� �I�7�m�[�}ϣϑ� ��A�s���߭���!� 3�i�Wߍ�{߱ߟ��� �������/��?�A� S�����y����� ���+��;�=�O��� s������������� 'K9o]�� ������5 #Yk߃��Q ����///U/ C/y/�/�/�/m/�/�/ �/�/?-???Q??u? c?�?�?�?�?�?�?�? OO'O)O;OqO_O�O �O�O�O�O�O�O__ 7_%_[_I__m_�_�_ �_�_�_�_o�'o9o �_o{oio�o�o�o�o �o�o�o/A�oe Su������ ���=�+�a�O�q� ��������ߏ͏�� ��'�]�K���o��� ��ɟ��ٟ���#�� G�5�k�Y�{���Ko�� ˯ݯ�����1��A� g�U���y�����ӿ� ��	���-��Q�c�u� ��Aϗϙϫ������ ��)��M�;�]߃�q� �ߕ��߹�������� �I�7�m�[���� �����������3�E� �]�o���������� ������-Se w5��������   �-�$TB�JOP_GRP �3����  ?�	hdEL�S�� ��`L� ��h X�0&���� @d	� �D�� �C�C�Y�xd�/?fff%�>��RD��@�@e-!B   A�dO/��x�/�/�%>���)!�?����"�33B; �?/�/c/u/�?%>��=$�9¹"���!� =!A���/p?� #@�6B�ffC�?�?�?>�%/5C�/ ^0@N0�1Y2�$�?w?�:�G�??OMJ333<��[C���3^@���"pOp�OO�?�HL���O�HY��>�@iB @��@N0yO_�O7W -_c7U_?_M_{_�_�_ A_�_�_�_�_o<oo �_[ouo_omo�o�o�C�N0 ��e	�V3.00jom9b7i*p�i%0w D��� E5� E߈` E�Kp�H� F\ F� FJpFL� F�cD Fz  F��^ F�� F��_p�` F�� F�. F�gp��� F�F@rE��pjp�� F��pG| G/ȿ GM G�pG߃� G��p�"� G�pG�n G�ͳpۺ G�q�� H� Hg) H�p�A<��KRP^1�aj#T�'�+�?�pa?_?� ��}������Ǐُ��� �!�3�E�W�i�{��� ����ß՟����� /�A�S�e�w������� ��ѯ�����+�=� O�a�s���������Ϳ ߿���'�9�K�]� oρϓϥϷ������� ���#�5�G�Y�k�}ߠ�ߡ߳�ahe��f�12345678�����[�=uEZ� �E�� F$ �F*�F�� F��3�h F.��� G� Gd� G2�G1� G�?h�s*�Ghl {GvK��� G:� %�7�I�[�m�=�p��M>� ?�C��	����?�4�F�=CPPACTSW��|S\�IR ���]  CH�_�SPEED 堋� ���  ��DY�_CFGG ���z����z����D%B���@�^09� "V�_CUR_�IDXl���V_E�XT_ENB  �w_HI�ST_BU 3�~Sd � �F��T�k �\�U`�d�h�l�TV� t�x�|�Tff� ������U��������T^4�������E����w����D�a����6� ��U��������U��������TZ0�������� ��0�����
P������������ *��$��(��,��s"��4�����<������������L�8�������%�1=IU�amy������R��)858A8UM8Y8e8q8U}8�8�8�8��8�6_MAX�_AN� n�_S�PD��o  ��xa:�o�pB�]O�UNUM��� s	
�WOUT {3�o	 
 55 GjAoSo�owo�o �o�o�o�o�o&�+=Oxa�ZERO��P�\�ESTPA�RSl���Ra�HR��pABLE 1�)kI�[@� �gwgxgx�'��gw�
gxgx�&�Qgx�gxgx2�rRDI�y�����/���O������͏ߏH���rS��w a� ğ֟�����0�B� T�f�x���������ү ������]����x �wMJ�\�n���,�>��P�b�t����rA�a U��#�  ����r�����ٱ�1�@a�IMEBF_�TT�qҵ�	o�VE�R�� ��l�R {1�)k 8�_����� ��f��� ���������"�4�F� X�j�|ߎߠ߲����� ������0�B��f� x������������� ��,�>�P�b�t��� ������������ (:�^p�������F���g�q@�erPMI_CH�ANx� e FDOBGLV�05�V�FETHERADW ?�U�����0�:e�4:�75:d8:f8� �9�fa�feb�R#`��!�Z�!�/�YISN�MASK�c�255.W%e3U/�g/y/e3rPOOLOFS_DI�p�z�u�ORQCTRL ��)k�����/��T �/?-???Q?c?u?�? �?�?�?�?�?�?OO )O;OKL�/nO]O�O��PE_DETAI�o�&yqPGL_C/ONFI�P�*�:����/cell�/$CID$/grp1�O__0_B_�T_����M/$F�P$/svgun [_�_�_�_�_`[�o o'o9oKo]o�_�o�o �o�o�o�ojo�o# 5GY�o�o��� ���x��1�C� U�g����������ӏ���k�}��'�9�K��]�o���ﱃO����� ��ޟ���&�8�� \�n���������E�گ ����"�4�F�կj� |�������ĿS���� ��0�B�ѿf�xϊ� �Ϯ�����a����� ,�>�P���t߆ߘߪ� ����]�����(�:� L�^��߂������ ��k� ��$�6�H�Z� ��~���������������@�User� View �I}�}1234567890-?Qc`u}�C���	2	z���'9��3��������@/�4 v;/M/_/q/�/�/��/�5*/�/??%? 7?I?�/j?�6�/�? �?�?�?�?�?\?O�7�?WOiO{O�O�O�OO�O�8FO__/_�A_S_e_�O�_�R �lCamera
_�_�_�_oo%o�E�_Ooaosn �o�o�o�o�o�o�)  �V�	�_7I[ m�8o���$���!�3�E�W�~_� �Vu�����Ǐُ� ���!�3�E���i�{� ������ßj�|�))Z� �!�3�E�W�i���� ������կ����� /�֟|�{ȯ}����� ��ſ׿~�����j� C�U�g�yϋϝ�D��U �92�������/�A� �e�w߉��ϭ߿��� ������|�EI��S� e�w����T����� ��@��+�=�O�a�s� �|��I
��������� ��=Oa�������������9 k 2DVhz! ���i��
//P./@/R/�J	�U0� �/�/�/�/�/�/�? ?/?�S?e?w?�?�? �?T/f/�P�[Q?OO *O<ONO`O?�O�O�O �?�O�O�O__&_�? �U{�Or_�_�_�_�_ �_sO�_oo__8oJo \ono�o�o9_s%��)o �o�o&8�_\ n��o����� ��o�e�J�\�n� ������Kȏڏ�7� �"�4�F�X�j���e ^����ȟڟ���� ��4�F�X���|����� ��į֯}��e��m�"� 4�F�X�j�|�#����� Ŀ������0�B��  �qσ� �ϧϹ����������%�7�   �)��C>�)C���@28B+��]��D��M�l�D��'?������7hDw9�5ߏߡ߳����� ������1�C�U�g� y������������ 	��-�?�Q�c�u��� ������������ );M_q����9�  
�(  ��e�( 	  ���7%[ Ikm����t��
G� ̑� B/T/f/ٿ�/�/�/�/ �/�/�1/? ?2?y/ V?h?z?�?�?�?�/�? �?�???O.O@OROdO vO�?�O�O�OO�O�O __*_<_�O�Or_�_ �_�O�_�_�_�_oo [_8oJo\o�_�o�o�o �o�o�o!o�o"io FXj|���o�o ���A�0�B�T� f�x���������� ����,�>���b�t� ��͏����Ο���� K�]�:�L�^������� ����ʯܯ#� ��$� k�H�Z�l�~������ ƿؿ�1�� �2�D� V�hϯ����ϰ���	� ����
��.�@߇�d� v߈��Ϭ߾������� �M�*�<�N��r�����������@ A������������ ��(frh:�\tpgl\ro�bots\m90�0ibY�_7\�f.xml������� �������� $1	�� I�dummy Um�r�����@��&=�- Rdv����� ��///)/N/`/ r/�/�/�/�/�/�/�/ ??+/%?J?\?n?�? �?�?�?�?�?�?�?O '?!OFOXOjO|O�O�O �O�O�O�O�O_#O_ B_T_f_x_�_�_�_�_ �_�_�_o_o>oPo boto�o�o�o�o�o�o��o~8�n� ���C�<< A� ?�{YQ s������� ��'�U�;�]���q����������ۏ	����(�$TPGL�_OUTPUT s�!�!�4�� I�^�����n/�FSD���+?���+�D�pb� ������ҟ����� ,�>�P�b�t�������@��ί���9p���2345678901!�3�E�W�i�{�����
*nos�elect*3�D�3VS���[����:�Q��� hkB����Ƹ?�/hB�µ����� �?�QB �����z�����XOB4� ��.�@�R�d�vψ� ��'ϳ������������}�8�J�\�n߀� �*߶���������� ���F�X�j�|��&� �������������� B�T�f�x�����4��� ��������(P bt��0B�� �(�6^p ���>��� / /$/��Z/l/~/�/ �/�/L/�/�/�/? ?x2?��9p$$�� �t7b?�?�?�?�?�? �? O�?$OOHO:OlO ^O�O�O�O�O�O�O�O �O __D_6_h_Z_�_}4q�_�_�_�_�_ o�m@;5oGoAz ( 	 �_|ojo �o�o�o�o�o�o�o�o B0fT�x� ������,�� P�>�`�b�t�����Ώ���  <<�_��N��<�N� (�r�����ǟa� ӟ��ן�3�E���I� {��g���ï����� W��/�ɯ�e�w�Q� ������������� +��7�aϿ�ѿ�ϩ� Cϱ��Ϲ����'߅� K�]���Iߓ�m���� ��9�������G�Y� 3�}����w�����q� ������C���+�y� ��%�����������U� g�-?��KuOa ������) ;_q�Y�A ����/%/�/ [/m//�/�/}/�/�/ 7/I/?!?�/)?W?1? C?�?�?�/�?�?o?�?�O�?�?AOSO�)�WGL1.XML�o�M�$TPOF?F_LIM �`����FNw_SV�@  d��JP_MON ����D`�`2�ISTRTC�HK �ⅰF��_�BVTCOMP�AT�HOQ�FVWV_AR ��MrX.�D &_ �_`��B�A_DEFPROG %Y�%	S012S�SW01�_�L_D?ISPLAY�@^��RINST_MSwK  l �Z?INUSERE_�T�LCKNlkQUI�CKMENro�TS7CRE�`�PR?tpsc�TNaЬ`�i�B�`_�iST�CZ�E�QRACE_�CFG ��I�rT�P	�T
?���BsHNL 3��Z1qy[ �Rew �������zuITEM 3�Q{� �%$123?456789�P:�B�  =<B�h�z���  !�����PL�Տ�S6���Z�� ,���B���Ə��ꏪ� �����f�V�h�z��� ���n�����
�ʯ .�@�R�̯v�"�H�Z� ��f�������ؿ<� ���r�ϖ���q�̿ ������&���JϜ� %߀�@ߤ�P�v߈��� ���"�4߮�X��*� <��`�������l�� �����T���x��S� ��n���������,� >�b�"��2X�� �������:� �B���D ����6�Zl ~/P/�t/�/��/ / /�/D/?h/(?:? �/P?�/?�?�/�?? �?�? Od?O�?�?�? &O�?|O�O�OO�O<O NO`O�O�O�OV_h_�O t_�O_�_&_�_J_
o o�_2o�_�_o8q�`�Sq��j�g   ��j )q�o�Y
 �o�o�2�jUD1:\�?|���aR_GR�P 1�%�� 	 @!p��{��������~� �+�9��q?c�N���r�?�  ������ ԏ����
�,�.� @�v�d����������П��	Re,�>� �j����|�����¯ �&��J�3�n�W��� ���x�����ҿ���� ���*�P�>�t�b� �φϼϪ����H��� זaSCB 2��k e�b�t߆߀�ߪ߼������ߊlU�TORIAL ἠk&=�gV_C�ONFIG ���m$q�o"��L�OUTPUT ��i���������� �"�4�F�X�j�|��� �������������� "4FXj|�� ������0 BTfx���� ���//,/>/P/ b/t/�/�/�/�/�/� �/??(?:?L?^?p? �?�?�?�?�?�/�? O O$O6OHOZOlO~O�O �O�O�O�?�O�O_ _ 2_D_V_h_z_�_�_�_ �_�_�O�_
oo.o@o Rodovo�o�o�o�o�o �_�o*<N` r������o� ��&�8�J�\�n��� ������ȏڏv���� �*�<�N�`�r����� ����̟ޟ���&� 8�J�\�n��������� ȯگ����"�4�F� X�j�|�������Ŀֿ �����0�B�T�f� xϊϜϮ��������� ��,�>�P�b�t߆� �ߪ߼��������� (�:�L�^�p���� �������� ��$�6� H�Z�l�~��������� ������� 2DV hz������ �	.@Rdv �������/ */</N/`/r/�/�/��/�/�/�/�/?����!?3?1? ^?��?�?�?�?�?�? �? OO$O6OHOZO/ ~O�O�O�O�O�O�O�O _ _2_D_V_h_yO�_ �_�_�_�_�_�_
oo .o@oRodou_�o�o�o �o�o�o�o*< N`qo����� ����&�8�J�\� n�������ȏڏ� ���"�4�F�X�j�{� ������ğ֟���� �0�B�T�f�w����� ����ү�����,� >�P�b�t��������� ο����(�:�L� ^�pρ��Ϧϸ����� �� ��$�6�H�Z�l��{��$TX_SCREEN 2�55�0�}�HTTP://172.19.���13 F�x�:��H��4�UUЅ�$�{���:���������������h�ttp�� ' �4  ���Ш:��Q�� ��F �WS#1 �z��p�� ��� }��12:8080�������� ��^�' �%�WTC0�4�F�8J�\�^��/DATA.HT�M?D=20&S�=0&I=1&G�OTO=GO ������   1� set var� ��[3].$D�ESTINATI�ON = '��=	�� FLT����9#A��� }�{ߓ� ������������~� ��-?Qcu��� ����� ;�_q���� 0�T//%/7/I/ [/���/�/�/�/�/ �/b/?�/3?E?W?i?�{?�??�?�$UA�LRM_MSG �?��� �  ��?~�Wro�ng Path �Number�<I�nvalid S�election��;%EOp2A,De�d�5%EArgu�ment�<Tu�rn Table�/TrunPADo}s�AWaiti@�For Main�tenance A1@@�?�;�O�O_��7�A BGLo�gic Not �Runn�@UAp�p1)_;Z2I_;Z3i_;Z4�_;V_�O�_��_o�_/o�@Vis�PBystem�RI�n Auto Mo!oo�owo�o�o�o �o�o�o�o&J= nas����� ����F�9�j�]� ������ď���ۏ� ��0�#�5�f�Y���}�ட������:Ca�pwe6�QCom�plete�8W�eld� Tim�eoutGTi�p Dress �W	�FaultH�� Chang�eS��ater �Sav���Read�y�7E�At�@x�imumN�8J%�ntroll��T�ZGE�Mot�@�[�>�QStoppZBC�}D��quest���1�yILow��e�Magazine�R9PJ��U�I�z[�e�Remo���OpenZF"P��S�till����Cl�os����չFixj�����ڶ �ɟInstaР�Stef�0��4�����%�Dum�traXHAA�ű���#�Έ�Adv�A������Gun �Is�RFully���7Sp�P%�p�t!х�O��Tem���[E�n�mand62�E�ffm����K-Lif��Pr�ox��5F�O�Inocreaذ A���TD��E�\�surĻ@��i5C����ax�~E��'�J�i3��AC�heckS�AAMo�v�A�~�E�1��E� Empt��e����֟����� ��/�"�4�e�X���|� ������������+���%BID ToomlOղ LJ I1.�b
2pb
3�b
4�b@��j��`����@aH�� ���ab.bN�eW`N,�p��������Ni�E�ne�m Err�o����C�P�@G�,�8�24V{HC ID=15 Wi@�MUnlatchXZA��!<>�*L�% ��f(�Q�'���,�(`'�C��sm�! th�e GO��Cur�rr@LOut o'f Rk��3M(��ir��R=�@f(Unknown�A�@4A #�?�?�?�?OO�ODO7OhO��Flo�wDr��M�PDeconect��O�ĜA��GLdժ�FDS�!Home� - PhysiWcal0�p`��A=n�PElemI1'Pxe|G�@Bunk��wis Q�ty.���f�����AU	Qejx�E��E]Feedٸ\$RMcan	Qb��djuN`�qOVO�_�:�N R  Vali	d�\`4�_
o�_.o�!o3odowJRivFs#un�@�1��K��`�c�O�ťj���dps �F4��eCycJ���c	ԩ����� _Åc1Q�@VogZ �~�����	� �-� �2�Q�V���z�૏��ϏtMSe�aѡM�8�SCA )U���P��/eP�|$�Purm�G1��uccK�f�Co�ӏ��w�����̟ ������&��J�=� n�a�s�����ȯ��� ߯���F�9�j�]� ������Ŀ���ۿ� ��0�#�5�f�Yϊ�}� �ϡϳ��������,� �P�C�U߆�yߪߝ� ���������(��L� ?�p�c�u������ ������$��H�;�l� _��������������� D7h[� �����
� .!3dW�{� ����/�*// N/A/S/�/w/�/�/�/ �/�/�/�/&??J?=?�n?a?s?�?vI�$U�ALRM_SEV  ����1�� � &�0�1�1�2 �3�?C�2L�7IO O?L�42O�2O�O�O��O�H�1ECFG ���5� �ve@�  A�Q   B�vd
 �?���59_K_]_ o_�_�_�_�_�_�_�_��W�AGRP 2���K 0vf	 ���?6��e���:��5����Ǫþ��@�#_.c�HOo�?UI�_BBL_NOT�E ��JT��l���0����@�bDEFPR�OG ?%�; �(%CC_AUT01_OLDvo�5%�b
�o@+ dO�s��������fFKEYD?ATA 1��9/`�p �G�6 �g�y�P��������,(�����4([ INST ]���  OOK T��?�΀unTchsup@�B� utW������[EDCM�D�ß&�RE��FOğǟ����:�!� ^�p�W���{���ʯ����կ�$� ���/frh/gu�i/whitehome.png%�`c�u��������<�instN�޿����&ϵ�  =�lookͲT�[�m�ϑ����2�D�sgtch2Q�������%�7���1��l�~ߐߢߴ����<�edcmd�[�����%�7�B�/arwrg̿s�� ����J��������  �2�D���h�z����� ����Q�����
. @��dv���� �_�*<N �r�����[ �//&/8/J/\/3� a/�/�/�/�/�/�/� ??*?<?N?`?�/�? �?�?�?�?�?m?�?O &O8OJO\OnO�?�O�O �O�O�O�O{O_"_4_ F_X_j_�O|_�_�_�_ �_�_�_�_o0oBoTo foxoo�o�o�o�o�o �o�o,>Pbt ������� �(�:�L�^�p���� ����ʏ܏� �����6�H�Z�l�~���+����6���ן� 4�ş�$�3�,
�O���POINT �97X��� 6OO�K����	�ONF �hup���� CH�OICE]ܯޮTOUCHUP� 	�4�X�?�|�c����� ��ֿ������0�ϠT�f�Mϊ�i+��w�hitehome�c�����������poinb�N�`�r߄����I�i/look >�@�������� ��conf>�H�M�_��q����6�hoic���������#�&�=��toucɠ��@a�s�����������arwrg=����� +"�Oas� ��8��� '9�]o��� �F���/#/5/ �Y/k/}/�/�/�/�/ T/�/�/??1?C?�/ g?y?�?�?�?�?��^? �?	OO-O?OQOX?uO �O�O�O�O�O^O�O_ _)_;_M___�O�_�_ �_�_�_�_l_oo%o 7oIo[o�_o�o�o�o �o�o�ozo!3E Wi�o����� �v��/�A�S�e� w��������я��� ���+�=�O�a�s�� ������͟ߟ���� '�9�K�]�o������@��ɯۯ�����0���������6�H�Z�2�|���h�, zϿ�r��ʿ�� � =�$�a�s�Zϗ�~ϻ� �ϴ������'��K� 2�o�Vߓߥߌ��߰� �����?#�5�G�Y�k� }����������� ���1�C�U�g�y��� �����������	�� -?Qcu��( �����; M_q��$�� ��//%/�I/[/ m//�/�/2/�/�/�/ �/?!?�/E?W?i?{? �?�?�?@?�?�?�?O O/O�?SOeOwO�O�O �O<O�O�O�O__+_ =_�a_s_�_�_�_�_ �O�_�_oo'o9oKo �_oo�o�o�o�o�oXo �o�o#5G�ok }�����f� ��1�C�U��y��� ������ӏb���	�� -�?�Q�c�򏇟���� ��ϟ�p���)�;� M�_��������˯ ݯ�~��%�7�I�[� m���������ǿٿ� z��!�3�E�W�i�{��RP���RP����ϸ��͢�������,��/���S�:� w߉�p߭ߔ������� ���+�=�$�a�H�� ��~��������� ��9� �]�o�N_���� ����������#5 GYk}��� ����1CU gy����� �	/�-/?/Q/c/u/ �//�/�/�/�/�/? �/)?;?M?_?q?�?�? $?�?�?�?�?OO�? 7OIO[OmOO�O O�O �O�O�O�O_!_�OE_ W_i_{_�_�_._�_�_ �_�_oo�_AoSoeo wo�o�o�o���o�o�o +2oOas� ���J���� '�9��]�o������� ��F�ۏ����#�5� G�֏k�}�������ş T������1�C�ҟ g�y���������ӯb� ��	��-�?�Q��u� ��������Ͽ^��� �)�;�M�_�ϕ� �Ϲ�����l���%� 7�I�[���ߑߣߵ���������`l��>�`����(� :��\�n�H�,Z��� R������������ A�S�:�w�^������� ��������+O 6s�l���� �o'9K]l� �������| /#/5/G/Y/k/��/ �/�/�/�/�/x/?? 1?C?U?g?y??�?�? �?�?�?�?�?O-O?O QOcOuOO�O�O�O�O �O�O_�O)_;_M___ q_�__�_�_�_�_�_ o�_%o7oIo[omoo �o o�o�o�o�o�o �o3EWi{� �������� A�S�e�w�������� я�����+���O� a�s�������8�͟ߟ ���'���K�]�o� ��������F�ۯ��� �#�5�įY�k�}��� ����B�׿����� 1�C�ҿg�yϋϝϯ� ��P�����	��-�?� ��c�u߇ߙ߽߫��� ^�����)�;�M��� q�������Z�����%�7�I�[�2�����2������������������,��3Wi P�t����� A(ew^ �������/  /=/O/.�s/�/�/�/ �/�/���/??'?9? K?]?�/�?�?�?�?�? �?j?�?O#O5OGOYO �?}O�O�O�O�O�O�O xO__1_C_U_g_�O �_�_�_�_�_�_t_	o o-o?oQocouoo�o �o�o�o�o�o�o) ;M_q ��� �����%�7�I� [�m�������Ǐُ �����!�3�E�W�i� {���d/��ß՟��� ��/�A�S�e�w��� ��*���ѯ����� ��=�O�a�s�����&� ��Ϳ߿���'϶� K�]�oρϓϥ�4��� �������#߲�G�Y� k�}ߏߡ߳�B����� ����1���U�g�y� ����>�������	� �-�?���c�u����� ����L�����) ;��_q��������L��������<N(,:/2/� ������!/3/ /W/>/{/�/t/�/�/ �/�/�/?�//??S? e?L?�?p?�?�?���? �?OO+O=OLaOsO �O�O�O�O�O\O�O_ _'_9_K_�Oo_�_�_ �_�_�_X_�_�_o#o 5oGoYo�_}o�o�o�o �o�ofo�o1C U�oy����� �t	��-�?�Q�c� ���������Ϗ�p� ��)�;�M�_�q� � ������˟ݟ�~�� %�7�I�[�m������� ��ǯٯ����?!�3� E�W�i�{�������ÿ տ���Ϛ�/�A�S� e�wω�ϭϿ����� ��ߖ�+�=�O�a�s� �ߗ�&߻�������� ��9�K�]�o��� "�����������#� ��G�Y�k�}�����0� ����������C Ugy���>� ��	-�Qc u���:����//)/;/��}�����f/@x/�-b/�/�/�&,�? �/�??�/7?I?0?m? T?�?�?�?�?�?�?�? �?!OOEOWO>O{ObO �O�O�O�O�O�O�O_ /_�S_e_w_�_�_�_ ��_�_�_oo+o=o �_aoso�o�o�o�oJo �o�o'9�o] o�����X� ��#�5�G��k�}� ������ŏT����� �1�C�U��y����� ����ӟb���	��-� ?�Q���u��������� ϯ�p���)�;�M� _��������˿ݿ l���%�7�I�[�m� D_�ϣϵ�������� �!�3�E�W�i�{�
� �߱��������߈�� /�A�S�e�w���� �����������+�=� O�a�s���������� ������'9K] o��"���� ��5GYk} ������/ /�C/U/g/y/�/�/ ,/�/�/�/�/	??�/ ??Q?c?u?�?�?�?���,;�������?�?�=�?O.OF,__O_�OjO�O �O�O�O�O__�O7_ _[_m_T_�_x_�_�_ �_�_�_o�_3oEo,o ioPo�o�o~��o�o�o �o,?ASew ���<���� �+��O�a�s����� ��8�͏ߏ���'� 9�ȏ]�o��������� F�۟����#�5�ğ Y�k�}�������ůT� �����1�C�үg� y���������P���� 	��-�?�Q��uχ� �ϫϽ���^����� )�;�M���q߃ߕߧ� �����ߴo��%�7� I�[�b������� ����z��!�3�E�W� i�������������� v�/ASew ������� +=Oas� �����/�'/ 9/K/]/o/�//�/�/ �/�/�/�/�/#?5?G? Y?k?}?�??�?�?�? �?�?O�?1OCOUOgO yO�OO�O�O�O�O�O�	__�$UI_I�NUSER  ����<Q?�  _ _�_MENHIST� 1�<U_  (KP���(/SOFTPA�RT/GENLI�NK?curre�nt=menup�age,153,�1  C�PSPO�T�Q�_�_�_ o�B)��_�^381,10
�R �Q4o^opo�o�o#o5i�P_S23>`  �_�o�o�o|�o5i2 NGE�a@�RVhz��B'!j37�Q0�a32�P T����E2��U�edit�RTIPDRES�g\�n���䒏�D-)�;�STY�LE01�q�p0R�BT�r���
���q/����ՀSSW�p93 Qr������G���@�Q����џ�����+� ��P�b� t�������9�ί�� ��(���L�^�p��� ������G�ܿ� �� $�6�ſZ�l�~ϐϢ� ��C�������� �2� D���h�zߌߞ߰��� ������
��.�@�R� U�v�������_� ����*�<�N���r� ������������m� &8J\���� ����i�" 4FXj���� ������/0/B/ T/f/x/{�/�/�/�/ �/�/�/?,?>?P?b? t??�?�?�?�?�?�? O�?(O:OLO^OpO�O O�O�O�O�O�O _�O _6_H_Z_l_~_�__ �_�_�_�_�_o��_ DoVohozo�o�o�_�o �o�o�o
�o@R dv���;�� ���*��N�`�r� ������7�̏ޏ��� �&�8�Ǐ\�n����� ����E�ڟ����"��4�k�$UI_P�ANEDATA �1����e��  	��}http:/�/172.19.���12:8080�/ cgi _h�eight=10�0&_devic�e=TP&_li�nes=3��columns=4���fon��4&_p�age=doub�1A�f)prsim��  }��4�F�X�j�|��� ) ������ؿ������� 2��V�h�Oό�sϰ���ϩ���f��� � ��}��/frh�/cgtp/TP�GL1.stm �m?_width=������2����Ѧy2���dual�� �� ���������+� ��O�6�s��l��� ���������'��K��]�D������ ��  ���xe����flex��'�-ߟ�3N�ʡZ�˥�t��3��k�hird$N��r��� ��s���& J1nU����@����"/�� h� F%g�bg/y/�/�/�/ �//�/X	??-??? Q?c?�/�?�?�?�?�? �?�?�?O�?;O"O_O qOXO�O|O�O�O>/P/ __%_7_I_[_�O_ �/�_�_�_�_�_�_o v_3ooWo>o{o�oto �o�o�o�o�o�o/ A(e�O�O��� ���H�+��_O� a�s��������͏�� ���'��K�]�D� ��h�������۟�� r�B�G�Y�k�}��� ����ů8������ 1�C���g�y�`����� ��ӿ����޿��?� Q�8�u�\ϙϫ��0� ������)�;ߎ�_� ү�ߕߧ߹������� V����7��[�m�T� ��x���������� !��E������P��� ����������)w� {���4FXj|� �������� 0TfM�q�����s������$�UI_POSTY�PE  ���� 	 ��H."QUICK�MEN  %+� H/L/_RESTORE 1����  ��*defa�ults�  I�NGLE�-P�RIM�/mme�nupage,9�61,1 ANG?E_S2330?�1?C?U?�)  5154?�?�?�?�?k8��?�?	OO-O?O  �NO`O�?�O�O�O�O �O�O�O_+_=_O_a_ _�_�_�_�_�_xO�_ �_�_p_9oKo]ooo�o $o�o�o�o�o�o�o�o #5GYkox� ������� C�U�g�y���.����� ӏ�������(��� L�u���������`�� ���)�̟M�_�q�x����O-SCREe �?j-u1�sc� u2֤3�֤4֤5֤6֤7r֤8֡��TAT!-�� y#��*US#ER����ϢT��أSks�q�4q�5q��6q�7q�8q� N�DO_CFG a�%+`�_� PD��S��No�neX"J�_INF�O 2�����w 0%���s��G� *�k�}�`ϡϳϖ��� �������1�C�&�g��N,�OFFSET' �%)�t�;� � D����������� $�Q�H�Z��^��� ���������� �2� |�z/~�l���
�����4�Ʊ�WORK ���6/��$u߾�UFRAM� ������RTOL_�ABRTe�}E�NB�wGRP �2Ϫ)v!Cz  A������� �"4FXyd �U����MSK � �����Nb�%���%N���_'EVN� ����v��3Ж�
 h���UEV� !�td:\event_user\�FI C7N/��>�F���B SPG!L'sp�otweld~-!�C6:\EVE�Ng�POTWELQD~/�/>��!� ]/?P?�'�	???-? �?�?c?u?�?�?O�? �?�?ZOO~O)O;OqO �O�O�O�O�O�O2_!_ V___�_7_�_�_m_�_�_�_o�_�Z&Wf��3�T���8o�o�o no�o�o�o�o �o�o#5YkF ��|�������1�C��T�y�����$VALD_CP�C 3Җ� qg�Ώ�� K� Ρ8&��3�E��;�.�dl�i�f��h� 4���4���џ���� �+�=�O�^�p����� ����ͯܟ�$��� 9�K�Z�l�~������� ��ۿ���� �5�G� ޿h�z�����Y�¿�� �������C�U�d� vψϮϬϾ���^��� ��*�?�Q�`�r߄� �ߨ߽���������� &�'�M�_�n���� �����������%4� I[j�|�������� �����!0EW ix��B��� �//>S/e/t �����/��// /+?:/O?a?s?�/�/ �/�/�?�/�? ??H? 9O(O]OoO~?�?�?�? �?�?�O�OO O5_DO Y_k__�O�O�O�O}_ �O�_
__�_@_2ogo yo�_�_�_�_�_�_�o �oo*o?Nocu�o �o�o�o�o��o� &�JK�q����� ��ʏ���"�4� I�X�m��������ď ֏�����0�E�T� i�{���������f�ԯ ����,�>�S�b�w� ��������ί���� �(�:�O�^�sυϗ� ����ʿܿ�� ��$� 6�l�]�L߁ߓߢϴ� ����������#�2�D� Y�h�}��&������ �ߡ�
��.�@���d� V�������������� ���<�N�cr�� ����������� )8J1no�� ��� �%/4 FXm/|�/�/�� ���?/3?B/T/ i?x/�?�?�?�/�/�/ �?�??/O>?P?b?wO �?�O�O�?�?�?�?O _(O=_LO^Os_�O�_ �_�_�O�O�O _o$_ 9oH_Z_�_�opo�o�o �_�_�_�_o o"G Voho}�o��J�o �o�o
�.C�Rd ��z�����������)��$VAR�S_CONFIG� �e�L��  qH  *�  �0��CMR_GRP ;2�L�Ԉہ�	ـX�  %1�: SC130E�F2 *����0��d0�e��؈ۀ�53��؁?�  A@���p���*� "���)�8�J�w�p��r����A�������3���ܯ3�? B�����3� �����c�@��d�O� ��s��������9�ÿ ���N��rτ�Ќ ������ԟ���
� '�.�K���T߁�8ϥ� �����������#�5� |��k�V������ ����@����1��U��\�y���3�IA_W�ORK �L���v�ۆ,		�f�L�����G�P ����U���SION�TMOUT  �0�S��  ��_CFG ��Q�S<�V� FR:�\\DATA\��� �� M�CNLOG[  � UD1NEX�3�' B@ ����9����)� �� n6  ����)��֌#��  =���Z0�W�� tTRAINة"i 
�pZ^�Y�e�.x��L� (G�� ?��//(/:/p/^/ �/�/�/�/�/�/�/�/^��S_GE6�L�7�`3��
v�t�,':� RE9 �L�E.4�LEX54�L�ـ�1-e��VMPH?ASE  L�؃���8�RTD_FILTER 2�~� �����O'O9O KO]OoO�O�O�O�O)�  O�O�O	__-_?_Q_�c_u_�_3�SHIF�TMENU 1�^L�
 <g�%��_ ���_�_"o�_ oXo/oAo�oeowo�o �o�o�o�o�oB�	LIVE/S�NA��%vsf�liv�>T�> SETU��wrmenu��,����U6�L�) �W+MO6�>�	�<�KZD"��q?d<���P�$WAIT?DINEND؁|6���OK  ��Ȧ�
��SՏ��TI]M�� �G�� "���E�ԏ%��%����RELE�1U�2�؋�'�_ACCTjpT���_W� ���%�ITPATH��_	��RDIS�p֞�7$XSh��n���p��Z�;Ԧ�XVRh���L��$ZAB�C�1�n� ,�J�2]�9��>����d��VSPT q�L���d
�z���������T�D/CSCH����C�M�ڸ�IPg��n�I�Q�c�u�N��MPCF_G 1왫 0B-��� �ϲ��ω���-���pB�G�E߀���@  ?��˺:��;Pߟ:9��d��:��9��aY�����dоD�1��ĐbKC%O�,d04ѿ�?����g!�:����5˿Ǫ�Ͼ��P�b��;�Q�p�:6��bF�� F���8�Ԯ���5Ǭ�Z؁�9�,�J�4�q���E�ټ�����D��I&:
��:;��B���������':�:':�Р���=��� ��������&���������;���W�2߳��������P� �G�Y����(�6L�{ *L�T��x��� ��>8Jtn,� ��'l�ޤ��90��-�	$_CYLI�ND�1�� ��� ,(  * [/l-%�X/�/|/�/�- �/?>U/6? �/Z?A?S?�?�/�?�? �??�?�?}?2OOVO�=O�?�O�O,�2���!� ����O�� �_�C_�S_y_]T��QA�b_�_�O4_ �_0_oT_�_;o�_+"�SPHERE 2�;-��?�o@O�o�o �o�onOEo 2�?V �o�o�s��	� �?Q.��R�9�K���������Џ�ZZ� �ߖ