��   ��A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ����PMC_CF�G_T   �� $'NUM_�MSK  $�EXE_TYPE�CMEM_OPT�PN_CNFCI�F_CY:gSC�N_TIME �E RESET_PȂDo LJ �HECK_DSBLC �$DRA> AR�GINCSTOR�JDISPKNETF_MISCCw�4&DEV._ d 	7OC�'HARADD�SIZORACnBSLO[ODK�IOKOCCPY�C&l /  L ��-UUI�DXC�L. 7� 
�EQPLnHRAT�TRK�BUF| .��U�N_STATUS�CU  �MAX�8(I��SNP_�PA�  �{ � ANNE��� Os CTION�_�PU�  � $BAUD��NOISY�NV�T1�#2�#3�$7_PR�T4PC �DATA�CQUwEUE� PTHw$�MM_ �%B!RE�TRIESCAU�TO)!R[��B�G) � ��INF���' CLIMI� ^5AD_H _3H ��#�6�#�6�#�6�# s1� �#�4�#�4�#�4��"� �$$CLA�SS  �����1�����0V�ERS� �8  1N���FG0 �5A���&@GAB�����d��OF��,C�  �38GC@d $ ED�O���O�O�O�O�O __:_)_^_M_�_q_ �_�_�_�_�_�_oo 6o%oZoIo~omo�o�o �o�o�o�o�o2! VEzi���� ��
��.��R�A� v�e����������я ���*��N�=�r�a� ��������ޟ͟�� &��J�9�n�]����� ����گɯ���"�� F�5�j�Y���}����� ֿſ�����B�1� f�Uϊ�yϮϝ����� �����	�>�-�b�Q� ��uߪߙ��߽����� ��:�)�^�M��q� ������������ 6�%�Z�I�~�m����� ����������2! VEzi���� ��
�.RA ve������ /�*//N/=/r/a/|v,,CIF 3�KWP EDFQHU@m�/|/�/?
??.? W?R?d?v?�?�?�?�? �?�?�?O/O*O<ONO wOrO�O�O�O�O�O�O ___&_O_J_\_n_ �_�_�_�_�_�_�_�_ 'o"o4oFooojo|o�o �o�o�o�o�o�o GBTf���� ������,�>� g�b�t���������Ώ �����?�:�L�^� ��������ϟʟܟ�����)TYPE �3�+ (�#R�!d'� �� #�"���ů� ���� ܯ�'�9��#S�NP_PARAM' �+����  '� ���@� ۠��"���� Uh��!ιݺ