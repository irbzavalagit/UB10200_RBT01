��   �E�A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ����DCSS_C�PC_T  �4 $COMM�ENT $�ENABLE � $MODJG�RP_NUMKL�\  $U�FRM\] _VT�X M �   �$Y�Z1K �$Z2�STOP�_TYPKDSB�IO�IDXKE�NBL_CALM�D�USE_PR�EDIC? �EL�AY_TIMJS�PEED_CTR�LKOVR_LI�M? p D� L�0��UTOOi��O^�4&S. � 8J\TC�u
!���0\� jY�0  � �C�HG_SIZ��$AP!�E�D�IS�]$!�C�_+{#s%O#J�p 	]$Jd#� �&s"�"{#p�)�$�'�_SE_EXPAN#N��iGSTAT/� DFP_BASE $0�K$4!� .6_V�7>H73hJ- ǌ }�\AX�S\UP�LW��7���a7r �< w?�?�?��?��?�//	7ELE}M/ T �&B.2NO�G]@%CN�HA�DF#� $DATA)he0 � PJ�@ �3 
&P5� �� 1U*n   _VSiSZbRj0RjR(�VyT(�R%S�{TROBOT�X�SARo�U�V$C�UR_��RjSE�TU4"	 }$d P_MGN�INP_ASSe# �PB!� `CiH�77`�e�.fXc1�CO�NFIG_CHK�`E_PO* }dSH�RST�gM^#/eOTHERRBT�j#_G]�R�dTv �k|u�dVALD_7hX�e�4hT1r
0R� HLHt� 0  lpt<NerRFYhH�~t�5�1� ��W\�_A$R� �T;PH/ (G%�Q�Q�Q3?wB;OX/ 8�@F! �F!�G �r��su�UIRi@  �,�F�pER%@3� $�p �l�_Sf�A�Z}N/ 0 IbF(@�p��Z_�0 _�0?wu0  �@�QWyv	*��~4��$$CL`  ����!���Q���Q�VERSI�ON� � 1N�$' �3 ?�Q  �Cell �Perimeteqr��J��� "��(��������1� E����������� E9�������ـ EӅ ����  yd��Cz  2����Z���u�m�anent Space 1`���Ǜ ����ğů������ +�=�O�a�s�2d��� ����ͯ�����'� 9�K�M�o�}�3hϛ� ����ѿ����
��+� =�O�Q�s�}�4lߟ� ������������/� A�S�U�w�}�5p�� �������� ��!�3� E�W�Y�{�}�6t��� ��������%�7� I�[�]�}�7x�� ������); M_a�}�8|� ����//-? Qce/�}�9�/� ��/��/?"?1/C/�U/g/i?�%Monitoring}� �/�/|?�/�?OO.? @?R?x?v?�?�<���? �?�O�?__*_9OKO ]OoOq_�O�5�ϿO�O �_�O
oo.o=_O_a_ s_uo�_�5���_�_�o �_ 2AoSoeowo y�o�5���o�o��o �$�6�EWi{}� ��5������� (�:�I�[�m������ �5�Ϗ�����,� >�M�_�q��������5 �ӟ���	��0�B� Q�c�u��������5�/ ׯ����"�4�F�U� g�y����ϋ%����ۿ ���&�8�J�Y�k� }Ϗϑ߳�������� ���4�F�U�g�yߋ� �߯����������� 0�B���c�u���� ����������	> P_�q���������� Y��%:L[ m������ �/!6/H/Z/i{ ���/��/��/  ?//D?V?e/w/�/�/ �/�?�/�?�/?O+? @OROdOs?�?�?=O�O �?�O�?OO*_9ON_ `_oO�O�O�O�O�O�_ �_�O_&o5_Jo\ono }_�_�_�_�o�_�o�_ oCo4#Xjyo�o �o�o�o�o��	 0�?T�f����� �ҏ�����я;� -�b�t�������͏ˏ�݊�$DCSS_CSC 3����Q � P����<�މd �m�0���T���x�ٯ �����ү3���W�� {�>���b���տ���� ����A��e�w�:� ��^Ͽς��Ϧ���� ��=� �a�$߅�Hߩ� l����ߢ����'��� K��o�2���h����������GRP ;3�� ����	ԟU�@�y�d����� ��������	��? *cN�r��� ���M8 q\������ /�/7/"/[/F// j/�/�/�/�/�/�/? �/?E?0?i?T?�?�? �?|?�?�?�?�?	O/O OSO>OwO�O�OfO�O �O�O�O_�O_=_(_ a_s_�_P_�_�_�_�_��_�_o'ooKo�_�GSTAT 3���M��< ���9�����뺸/{�`�:�:���]�;nS:����`��C΍Đ���Dg�f��:`<��e>���q&��4��p3�EI?�  �a���`4��ZC	�o����`  ����e�	�>���?ho}���}?Z�֑��i��g`B_��`D~9�z���7?q"<:�ʙ�z��</������i���5BC�lA��cy:����?#�?��Jw�M�`������5_C�'��Đ�pD����y>��Z�`�����?�p�p�;5��h�����?�b��o �o�ow��>�P���2� |���h���ď҉�i�a /i�-ky�0��zU�p~t�"p �i�ÇҗD>�lD�.�"�D���X� ���ʟܟ��,���\� n���z���~���گ� �0��D��L�2�@�Rp�Vp�Zp^p�
&|h6t�B�d�οx� ֿ�����L�Ư|� �������Ϟϰ���߾^��7����`������69���6Χj�����6��I2�C����ďfDk�>�n��p����c^y3��x�bsоo��b:�$���Z���>�V%?h�x����?Zߊ��bʆ����P�Bn�D}���^�o�?s�6���5�86��*�2ц���`�C��w;����^�6���,���a����������6���C��}V�xD�!��z</�rѷ8D��n����06�ֿ���K�aF�(�:� L���������� ��� �V�h��Pϒ�dϊ�������߲߈�Ë��D?�D}�#����J��R�f x��B��
<� @,v�~����������1�����6�G6�ܩ����������� � /j//r/�/�/�/ �/�/b?*?\6?`? :?L?�?�?����X� j�|ߎ��������� ����0�B�T�f�x� ���?�?��?|_�_h_ �_�_�_�_�_��/�/ 6o�/>oloRoDOVO( ^o�o�oXo�o 8 V<�_���_�� ���(�olR�� Z���n� /2/D/z��� ����<�"�4�V��� ���Ɵ�ҟ��֟� 2�D�*_<_N_�?OO *O�o�o`OrO�O�O�O �O�O�O�O__&_h� z�\_&��*��N�`� :�lϖ�0�n�����h� ��������o��� ���ώ߼ߢ������� ~�4�F�x�j�|�V�h� �����������$� 
���Ώ���8���L� ���������� ��P b��n�r��� ƿؿ꿐�����Ư4� F���� �2�D�V�h� z�������¿�� ��/�/�/�/�/�/? 2?��
,n?v?�? �?|�`ߖ?�?"O�? *OXO>OpO�OtO?�O �O?__�O_N_`_ V?�O�_�O�_�_�_X� j�|��_�_>o�_Foto Zolo�o�o6_�o�o0_ 
4 j|b/t/ �/,>Pb�?�?� �����//(/ :/L/^/���/^P� b�<�����r���Οh_ �o�o
��o�@�&�� *��?2�T���,�Ư�� گ�*����l�~��� ������������@� &�T�.�\�B��_oo N�p��τ������� *�X�ҿ�ߚ�̿���� �߼������"�� ���l�~�4�F�X� j�|�������ď֏� ��<�N�0��������� "4@j�B�d� �<߮����� ��Z�b�v� ��R//L>/P/ */</�/�/���/� �/�/�/�Ϣϴ��/? v? ?~?�?�?�?�?�? n/$O6Oh/BOlOFOXO �O�O������d�v�� ���������� *�<�N�`�r������O �O���O�o�oto�o�o �o�o�/�? OB�? Jx^P_b_4j� �d�,��D�b�H� �o�����oڏ�Ə؏ "�4�*x�^���f��� z�,?>?P?������� �H�.�@�b���
��� ү�ޯ����>�P��B��$DCSS_�JPC 3B��Q ( D?`���������� ��ݿ��������� [�*�i�Nϣ�r��ϖ� �Ϻ����3���i� 8�J�\߱߀��ߤ��� �����A��"�w�F� X�j��������� +���O��0�r���f� x�����������9 ],�P�t� ����#�1 k:�^���� ���1/ //$/y/ H/�/l/�/�/�/�/	? �/�/??? ?2?�?V? �?z?�?�?�?�?O�? �?:O_O.O@O�OdOvO �O�O�O_�O%_�OI_ _m_<_N_�_r_�_�_��_�_�_��j�Ss��w�L�_Woo{o��d Fo�ojo�o�o�o�o �o3�oW{BT f������� A��e�,���P���t� ��������Ώ���O� �s�:���^�����ߟ ���ʟ'�� ��[� ��H���l�ɯ���� �د5���Y� �g�D� ��h�z�������¿� �C�
�g�.ϋ�Rϯ� v��ϚϬϾ��-��� Q��u�<ߙ�`߽߄� �ߨ�������M�� &�8�J��n������ �����7���[�"�� F�X�j����������� !��Ei0�T �x������ �Sw>�b�����/�(dMO�DEL 35k�x	Dres�spack/
 �<�j$�x �C/� ��  �*  . �  CH�'f/x$9*�'Ë!4� z�$�$
�c(z!�� Q/ ��/�/D??-?z?Q? c?u?�?�?�?�?�?�? .OOO)OvOMO_O�_SSW1�O^,�I�y#�%� ��8���!C�w!���X�Cu�Dg/5	�Ox$���&���V%�e2l�Dd���UƞBQÎk�_�O��ٽ�������C���B}խ�w�(V_�h_��J����Dd�������C>6�D|�鷒_x$��Ip����MC%�����DpC�C���O�O�O|Oo (ouoLo^o�o�o�o�o �o�o�o�J��M�o |�oew���� ��0���+�=�O� a�������䏻�͏ߏ ���b�9�K���3 Es����m�۟�:� �#�p�G�Y���}��� ���ůׯ$����Z� 1�C�U���y���ؿ�� ��ϩ���͟���� Q�cϰχϙ��Ͻ��� ������d�;�Mߚ� q߃ߕߧ߹������ �N�%�7�I�Ϩ�C� q��Y�����&���� \�3�E�W�i�{����� ��������/ A�ew���� ������f=O �s�����/ �/P/'/9/�/]/o/ �/�/�/�/?�/�/:? ?#?5?�?/]?o? �?�?�?O�?�?OO 1OCO�OgOyO�O�O�O �O�O�O�OD__-_z_ Q_c_u_�_�_�_�?
o �?�_�_Ro)o;o�o_o qo�o�o�o�o�o�o <%7I[m� �������� !��_��oI�[�ȏ�� ����Տ���F��/� |�S�e����������� џ�0���f�=�O� a�������m������ ѯ>���'�9�K�]�o� �������ɿۿ��� �#�p�G�YϦ�}Ϗ� �ϳ�����$����Z� ���5�Gߴ�/ߝ߯� ������2�	��h�?� Q�c�u�������� �����)�;�M��� q�����k�}߫���* ��%rI[� �����&� \3E�i{�� ��/��F/���� 3/E//�/�/�/�/ �/?�/??+?=?O? �?s?�?�?�?�?�?�? �?OPO'O9O�O]OoO �OW/�O{/�O�O�O�O _^_5_G_�_k_}_�_ �_�_�_o�_�_Hoo 1oCoUogoyo�o�o�o �o�o�o�o�OV�O 1�u����
� ���R�)�;���_� q����������ݏ� <��%�r�I�[�m�����$DCSS_P�STAT ����ՑQ�   �����  ��(�-��Q�n��  x� ��֐֐������������Օ�֯�ƔSETUP 	ՙ'BȘ�����:� T�ϯx�g����������I�ƔT1SC 3i
-�����Cz�����)��CP S-�D�DNt� ��@�ϼ��ϝ���� ���:�L�^�-߂ߔ� cߥ����߫� ��$� ��H�Z�l�;���� �������� �2�� V�h�z�I��������� ������	.@d v���`ϵ�N� ��3EW&{ ��n����/ /�A/S/e/4/�/�/ �/|/�/�/�/�/?+? �/?a?s?B?�?�?�? �?�?�?O�?'O9OKO OoO�OPO�O�O�O� �O�O_�O5_G_Y_(_ }_�_�_p_�_�_�_�_ oo�_CoUogo6o�o �o�o~o�o�o�o�o -�oQcuD�� ������)�;� 
��q���R�����ˏ ������O7�I�[� ������r�ǟٟ�� ���!��E�W�i�8� ��������կ篶�ȯ �/���S�e�w�F��� ����������ֿ+� =��a�sυ�Tϩϻ� �Ϝ�������9�K� ]�,��ߓ��t����� �����#���G�Y�k� :���������� ��1� �U�g�y�H� ���������������� -?cu�V� �����; Mq��d߹� �d//%/�I/[/ m/</�/�/r/�/�/�/ �/?!?3??W?i?{? J?�?�?�?�?�?�?�? O/OAOOeOwO�OXO �O�O�O�O�O_�O�O =_O__s_�_�_f_�_ �_�_�oo'o�_Ko ]ooo>o�o�oto�o�o �o�o#5Yk }L������ ��1�C��g�y��� Z�����ӏ����	�؏ -�?�Q� �u�����h� ��ϟ៰���)��_ M�_��@�����v�˯ ݯﯾ��%�7��[� m��N�������ٿ� ��̿!�3�E��i�{� ��\ϱ��ϒϤ���� ��/�A�S�"�w߉ߛ� j߿����߲������=�O�a�0��$DC�SS_TCPMA�P  ������Q @� 8�8�8�T8���8�8�8�U8�	8�
8�8�U8�8�8�9�W  8�8�8�U8�8�8�8�8�8�8�8��8�8�8�8� �8�!8�"8�#8�$�8�%8�&8�'8�(�8�)8�*8�+8�,�8�-8�.8�/8�0�8�18�28�38�4�8�58�68�78�8�8�98�:8�;8�<�8�=8�>8�?8�@��UIRO 3.��������� ���� $6HZ l~�������7���7��[ m������ �/!/3/E/W/i/{/ �/�/<�/�/�/? ?/?A?S?e?w?�?�? �?�?�?�?�?OO�/ =O�/aOsO�O�O�O�O �O�O�O__'_9_K_ ]_o_�_�_�_0O�_{�UIZN 3��	 �����
oo .o4�o\ono�oCo�o �o�o�o�o�o�o4 FX'|��c� �����0�B�� f�x�G�������ҏ�� �����>�P�b�%� ������y�Ο��򟵟 �(�:�	�^�p���E� W���ʯ��� ���_~��UFRM S�����8;�h�z� 9����Կ���
� ���@�R�-�vψ�c� �Ͼϙ��������*� <�S�`�r�ߖߨ߃� ���߹�����8�J� %�n��[������ ������"�4�K�X�j� 	�����{��������� ��BT/x� e������ ,C�Pb��s ����//�:/ L/'/p/�/]/�/�/�/ �/�/�/?$?;2?Z? l?G?�?�?}?�?�?�? �?O�?2ODOOhOzO UO�O�O�O�O�O�O
_ _3?E?R_d__�_�_ u_�_�_�_�_o�_*o <oo`oroMo�o�o�o �o�o�o�o&=_J \�o��m��� ���"�4��E�j� |�W�������֏�Ï ��5B�T��x��� e�������џ���� ,�>��b�t�O����� ��ί௻����