��  9��A��*SYST�EM*��V9.3�0126 2/�12/2021 A X  ���`�FC_CON�FIG_T  � @ $DAT�A_NUM  �$DUMMY1�B F2MEBU�GB $OUTPOS4INRLB w4&GRP0�� $FC�Tp  	� M_D_TRQ� � �SCH>�HOL�D�RESTAR�T�COMPLE�TE�MAX_E�RR_MM  ��IM_]FC?ENB_CN� d �DIZCMP�	S[TR�WT
S�)�2���W ����P
�FCGA�IN�? _��PS�/t_C?�MP��GUNCLOS�DFLa �TLM?OD_RQS�2��D_KG?�F�� ���R4M5�M�v:1  L�7 TIM� 
��
$EX_IN�PU�9"gA&TM_OBSERV�d7 wP%c  � ~" 3 j#�FB0 D q$�!� �	SIGh��EXTRA_L�ON�(!�#REAN� 
$� T0x �� ���'�$MOVE�R= HI�%REF�_A� �DIST�_1D��2�$W?ELD_ON�$�|j �CDDSB�"�*M5t_Ic#�4Z �CUR�INIT?_PRS_D[5�6�T�)�!1?�3' �1ATM1�1� ` �EDL�y2�TgASK>)ED� �DPT?+E�d P�:KNE+@REPL�Ah 4�SG�ATC* �� %$ATUNq_l@�d CS1>�_�  d GTS�JCS2�Kz@� |@�#$V_A�(!� �RL_VAL_IB �@_Mg�@l@��C�A�B�D?�FCCR�[ V�BUNOV_�THRH��AOyK� �@ADJ_'Q
�CLU�DQQ T� �UP_@EDB_V TUvR TvP�@z@�sS�@)P�VVASV�T�WD*0�V�P2�TxB�BT�O�@w�BT2 �G�TV�1� }S*0x�:dqARTQ�A�fPdLI
RgAXImACy"qb?�1g@�B y"�A�ffA)M�Pv`	�n	fA+P�K�v`
 � �$OPN_4TC̐PA$�`�`AF��`�bRE��`1L)Ob�fH�A�apB� C�Ss#w�d2�oW�g2|2wep#z�up#v!�`ME�F�G1_  0~^`OK2_CL��B&@�0SRC_�TY�A�sWb R�E �x2�p 8`� �}�A�s�0PD
���:�yua ��!D�ITO�0� N�U�@U1H��`NES*Bq J�P� ��!?$MEA)@/B��$Ep4�pINFvq$.BOFS�s1����A4�xBv`u5 : E_M�s���؀�r�䄸p2i1�a�"IN�0cD)� #$EwQUI~ YPE�B1DP�qa�"$�`|��b
qBTJ�A�q G1E��j�p�t�`l�	E�WIT� �UFA!d �2�=Q�$LPARA�
7 F��!�bH�X SRYg ڀK��D�90PQ�bSHO�aWsܠsi��aRD�_AT�0�eR�S�E!QE FL�RP� �xAH�$NOM�OT�PCSW�bC{LR84PMTaA @R��p�Db�W&B� BAS?0�2���`8�@��*�SUB�u�/SCRNՓL���N�;EQZ�#��Z;1gc���AC�phcޢ?FLENSCKcߡ_CUSTO��m�a�DG5� d >P_HKY_�AaO$BU@��D-��IF�Q�PG= FI1O�so�ID�C�A�CH�֓!SGD�IAskPv`� e$AV��p�b �� pLAP����ɳ� ���ƶ�ӸI��� ���ӷT�� ��1ǵ�Ws´Wͷ\� ݴWs�j�f��w�À��f�-�W9��õ�3 ����ͷ��ݴ����� ���
��%���-���,9�[�PR�X���b�n� p�Bnԇ���IN�u�IN��IN��C�OUNT� CדP�ROG_NA#!90{@YCL��Ep<���DO_Ns�5I�C�TVV* SECTI>1*0�OV7ae VHE���bUN5��`Y����RE �����h�0�� CCCA90���V�LV��v�IAG_�HO�1���E��AMuP
SL��YEAB�8������DAY�������DS��E�'��!�'�;���;���D��K�⦷0l�l�PCTT9OKc��FRC��y�EsF@�RSCQp�CQ ��CQ��CQ������Q�������6�x�LOK�$��1b�5 �r���_DL�x��p��C+~	SOL� p@����x�U�0�� �0	m�`�aD���PDE�A;�8r=�P(�E�pM@��E�p)3(eB��q�� xA" !��!! Aa|�_������ /�-1��EA��;��
�QS��Lt��b��o!�� (� 1 �p��OS�1# ��#���2 L�d�r��^���a��ض�a��E�RING_R������� �������h1���� �&$�%�*��(6�0 Q&"9e""5u��@%2CP~O4NEWUPDApR0�c�⬰ ��@�SW�`�@��V G1����5
}�0���7	78�0@m�CP�"��0�5��5
�ps41� �� p�DEVIC���UE����q�SI�Z�� ��Am�MAI�Nn�xs8��DEBU������I5��LO����C@���a�2��� �_$WRDW-�O�(E����FF��E.��b�OO��pCLOS;DIB�TIPW됏TROKİ�E�QUـ�R��a�� ����VaQERgd}�VER_OFF�|�}Q�INH_M�DTS�T(QTUq���s�_SPE5�Qm�����:�T1pב�SPUSH�Wi�ѐ�VQ���S
oPNiSs�ִ�V5��US,h(a\úV��Af Yh(a�úV[�Af�h(aA4-k�a?h�h(a5-k�a?h�h(a6-kq?hx(a7-k:q?h:x(aA8-kgq?hgx(a9-k �q?h�x(b�2g�?i �x(b,m;mJl1Yl!��?iwl1�lQ�?i�l1�l��?i�l1�l��?i�c_A�فɳ؂T\�؁B݇B,iDJR����@�U�C��ORIGINALe�AEh�A�GTHT�rhZ��\��Ct ��W��DOsWN�U&P_WD-� �TP���C&P���BP|�#��STNDR�S�����e��b���OUCHMET	H&PR�Pu�2��� P5�R���Ь�Εr�9E/Q~�CMPx�ܕ ����ܘq�ΥJ�q����΢Ct�&!�������.�&�TS_W�AIoT�Qp WI<,�* BF_V�Ro�G_�_D |����EXC��SYNCfo�DZo8�DZT&�DIZG@G&�IcZG�V$�@ME3�D���AE7���J�Iv�cFY8��J�CHy00S2þX5�AC��4��,�S4�DI8�DIb��E.�n!�OP`BL_�@]㫷����®��F2á���AUꐷ#��|Q��F�ާ�WSTP��THK�0Pޔ��s��DO$�Om ��:�I ��:��QT�Sӽ�8�z���z�PLu��OK�MS�Q�THCsKNUPF�FIXt MI	�UTb��Ab��CR �SB�h�T�E˶�M��t�#�R�EVOt�$LI�ۖSTo@���Pr6R>��REE�����Ҹ�& ��I��H�OL��C��I_ "% �@_�F��A �t��Yd��d��d��f�cSV��8�P_���NGtBQP_X&�_�/��/�Zѓ@�Q�$X�!�Z���\5 <UPLUO�T;V`���EQG@O j������PATl�H~PS 7�0�2��C�xX�1����WR��_f0 	�ԑ'n�����VTMP��S��P�g0��sP�X�  �C�AM`�Q�AM�ANU�Q  ���3_�,�U5�RK�J��3c��b0RBA�CK�@��RUSE��1dCn NA>P�%
�,!WELD F�GU�N��$'�5PT���y&�_T��J� B��>�@\ +�G�Dc�#�Q��e�DEP�T�S�C=�SOFTY_"�0SFT�A\S #��_P��%%")��o��S�z@CELs!+�J0L� B%f$O% 
 �&�$�$B&�#<O%�
AWAY@'�"�O%�l��U5U�~�O 7���W�7�-2-�e S�_  �!L4�"�L0-�U��e PATHN6t6��� ���\�c8ƌ��2�Q v�Ydv���:��DK���D[�R0�AI��@ ���I��˰J�v�vO%A�@�^@0 fG�U\BO%�𭵱�0E ��ܕ���4���Q�E�ΖQ	4�a\!IO~�   $d�P��Ռ �PE_��a��G�O�O���� < $'�F2�r�R2aS��1 
9$ayP 
5���Y��1�  t 	6�AB*�$�P7��I�PUL�0"U���l�_z��R����_M�ݱM�U���x E�� DPP�q��B<R0�_CMD.b`��*f��+j+`FR0O�pe�|��  Pn{�LON }P�|�RE�  
w  �TWD��!� B$BZ�� 5���S���Bn H�A\20�4�TO�OcRG�մ�TEƲ8�b}�v0LOA��k决RSӲ� j ZR�ӡ�0w �U� CST퓎��ȴF��Lds��@�M�|r�S�����RETRY_FL���aHPϒ��sIS�f�G_G<�n�pCLB��IS����QSKPRs�s^s�� ����B�7MTN�:��3Gŝ1W"��NWR_ATX��H�����35��H�,WB��`��͖��ܕ�b4W�Ts�DIV��OR�Kk3TWP�T��W�_PSH�PP�ET� ��r�LO�$�X΀D� F[�18�k�l�W_2��8��%���MEM��R�><FSTMCR�t��E���0 ~t�Qyy�_�`��N�$ZR�p_FR!~��Rs@���P0��fr�B� !F8`���ހD���s�RE!�0j ��T��8t�C�b"�mD��HRg�GA< Rp�g�q%��悥ŕ�wU��Z�v�0OLL�aCՔ��:� ��#�ΡAXԦsi!������JOG_VsEL��P GN4�s ��x����Ѹ�#� =e M_R���q���K1��`S�Z �!'�U3GRn@V<$��TupL����1�pOO���E�RVED���aLSzpE��MOSI
a
ߴE��CϠ߲��t��ERR��@�WEIKGH��X��T�ƀ$�7�K�a�'�A�'�EX7`H1~aj�&�'�}� 3�t�ȝ�n��0-�xnsSXK6_F� �����ՠL�$��DZ\Y���OVS��I��#K7gЎ0F�#҂��7���@�;�PAR@ }P�k���:�D��@a|�i %R ���P��dr�1�e����0IT������� ��3CV]'�0PF��f����`�EXTRA��~d�f$R�D_HPDFLT�R�do�0gM�@5OVR�Q�ѧƘ�ȵ�1���GF��i Z_O�F�D� ��sDOSp�$�`��^!�xB��]  P �Z �A0E�C=D�������Ƹ�CU��EX���A�%NP$ANLp1!�V���V��2]�20��A�IM��� & � $ ���1��KN��ô��3���3��4��5��6���7��8��9��10a�_PT4����#b�`8��`��NWTc��' 8 �M U�c��4w�3w|B�RSADJDB( 0ࢦ�0b��2Q$� _P�qQ��UTO�)� �j �UR`#�_ �c��4b�,6����a$D�pV2�dpZ�� k`ՃѡZuDZ��DA�p��
���÷�3w1~2
~1�2�A�A ,f��0<�5*?C�䓄"�T#_��a'��0CC_R2�%"�O#�S��k � ��yP( 
U�N��UPDVGS*� `����&�BSR�V<
�ARCH@sf�CЅ�႐a$�1�3�a� b�&�dLW�%+�/�/�/?d� >�G�AC�%,  �G6��_���ROBOTg4'��h38�&��DI#��PP[��T�&�F���7�A�CT DGSL�@J��(QI{4̠R���$ZD*�C�EU�T䠠�4+ rCN��N2x�T���sBSL[��@BN0ptP0q�LAt�&���be0P-� ��{�R�L�NCL&� E�2��1#��I��'���8�g2�APNL�`V�����USR&�(SP��CUAVo�n�S��b��PMP��%��aK��`r�bT+QWӁ�WG�WNUfQ�`70AS�UU�PASMXfPER_�NAKU�ORN�T�A�U���TRID5X�RPfUN*�1T/RKRE�W�C<QaT�'�7fA	ak��IZ!�b+�
6Sh�'�T8Q S��To�_EB*eM�edGӡ�cMP,pMVR��AL�� �e80L�(p r�c�� �i*`xE�b<a��d�0aM�� y���bTQ����eBS�`ÿ���4 �0zIvz�0vu�1�x
D�U�Rvu)��wv Ёvu���w�]`�w�a0�vN2���wBK�v3S��v�ALW�{LWC�TMG�wN1��4aL~�T�x�[�IN[�P�Ay�w�+�1��2[�:�TH[��B�@���IAS4AX��AgRML�p�DId�P�?PCR�p��� 񄍐W(QTDITUP7�2���琱4�a�㐰��l��a<� S�� ��Q��Г�4(q���ṘHK�k�z�X�q�ӤPLM����CCUT��j�𐹘�LM� j�c�!���81S�6�KPCဗvx|����BSTM7� 4Q���Q�k�sחY  Ԙ�@����o��w�@���ĊԒƅLINK1���2�3�1���G��C�-�G�P;�P� E񄱑v���@v0 vwA�v�}��@|�f@|�0�y�p� ��*ŵk��+$ABNOM����,�qBNWsAV���$��V��LG� t��� 7� �7�x�A�vw~f�p�P�A���SFRCU�CHCLB_CO;$��DON��Ļ�±�PZ"7 ǳws,$MBKLSH��?NMMAVG��ɷ���VGC��WRF�V�$qSA�sTRY_� H�SLT�0�wB�#OU& T�B�Fs0b�BpM�Aח���rL���a�0THO��`���� ��S��.t 8��Fq�#`��s�a � � 
z��B{t�Gp-D�tP@�z�l"?� �CZ�P`X��W�5 � 94H�-ITE��!�. FIp��CUR |&C�0�#��B. �`wF��_S�0��;�Wf�Vg���ma�gg���P1�Q�e�b�p��DYNTQv0�գ�D_ Ӯ����N �gcSHOR�t��r��G��e�M�'LBSP ӌ�jPPv0U8P�NUP48�HKLW��UR�F����@P��**	FUB�t*tPE{PHK4�@��CTD6q��ЄPaE��r1�ENT�B��U����0N��D��6`B���Wf3yֵT�t���ILNO�P5 l" �(Sl"IGNR�PT�H�	4�1EL�YWLD� / wl � ABL��EWU4�Q�Ps���F��PT����V6�yR���0$SWiQ���aT�BUN�INFO[0 @��0�ˁ�7�`�2�_!S5 �� �0D: ���1FCPAR}A�  1 �k��CTRL2�'REEP����v�q�c`3MP�fc!INA_q�d !�2b"V4�!F�NC_MSK��OM_��rV @ࠡ�9`_ y�C�2$o���0� 20�0L�Oq�FC2� _4TW�a3��#r!��q�2��-!2 �o1HK2iQ��02$�87OKMSQ�-2�R� �cS_3H2,2OK_PDf1Z�.0X��9��s_L�4�0_PLq���uT~� "!S�A�@ 3 � $�1�&��sb�1t�h�6�A�5ZqdTB���AL��AUSTO�R� �1a3A<�;Dp@��(DbhLON ��bot` �PLOT�CF�24 � ?$XAXIS�О%�p�`NS�P�K�����js��<sDBOUNCE�3`qP�`U��� b{��#�3�"!&�-!�5  �q�Ama�NU����.z fdAyPafe�Q�USb�TWѰ$�����R��$SG�RE � �P 2W!$C�Q"� U)�##m���Ѱ$f`��}AѰ%$SIM&��Ѱ&$NW�NG�i'�pMI4�O�_��)p Az-��^R.$(�LY_^X /6 _("RE`1��E`2�rA ��3$�DE`42N�RM�C6� ;$ROH�Y�r�%�Ύ`COR`1؃HA1P�@�ԭcRAV㇑�_XU��hN�Q�eY��jY�eb{�pr�OF�b��RLFx�aM�O�B�C���A�%�cOPj�e[#�`O�q2}`�sR��cuzr� ��6�DI�ӒwIDt�L�OC� TLUs>N`|�x��tW�MVqql��4B4}`PR����uN��%$AF@�{��������Z��f�zrRDY��zro�`��}`5�I��`4T��.�ADr C��ip��gSTRȰ��EN�*��I�� 4����@���������N��p��@Up�$$Z|�14MID*,�2�1�`G�fA�.�$POPUPWI:��;���DW����BL�NK�4LN���qBȃ㼑}`H�`��PRCME��t�C��_��HDV�P��OL4`0 `�����`IT�I��X��7 ( ���SXF �pA1�Pz�2=�3�=�O�`BUF�a8 D 	$RBX��yP7�Pk��$X�=�Y=�Z=�W=�P
=�R=�D=���E�!�~�`9( $��p�ХQi�{�TOU3�Xԑ>�e�_BxY��AT����з�褙O�=�HI�B�B4_��1����;�� H�N��R?���G�~�a n���z�zs�rФA���>�"pù���t}`��S�a: |b�zq��{p�a���`CHG_Wcᙢ�s���P�P%�b�ET�FLUC棾�UR�CY_E��}`E�X�@ ;x /-$US�0R{`���TSK_�����C����EQ��NQ��#DG�q��w�I��}c? 6$O��j �8o���A0��8$W	�`��؍`�!�p�X_$�=�p�Y8�Z8�$�c����?4_VX_V��p�P0j�Y������Q �¢Ԫ֝���2�T�ãX1��< ��Y��Y<�׳�39 �� 1V5w����KEV�v��Cr>����:��REQ�������������o�kᤀ ?,]J<�Z���r�>�5�_�IePSK��`��p��"p=�IIU�;FB-!< X���J�F�sr�����쑀U�f1Z�jO|C�2�=�
T �$ASSO3���VS�ư�X �M:�~�S��� O_CWAu Ѳ�6�����Q�USapTKL ��XX ���Y�@��Β M_E���$p����DOUh�� 	 ��Tq.Ǡ� 0ɣ!	 SG1 H!�P_0\
Ǡ��L0~d�ǠAU�Ц2�3p`�R��F* ��RX P�N@��j � 	(1_BU	H���P;�CjhAFDn�1�P	�1�@ 	���R�E���sYP� 0SPE)�ulq 'SE�@6�0z��M(DECE�P�d�`NE�cc]�p/]���/PATxPx10j DTCT��PEPPM��p�="��"O02A�2��`U�N�-pT ASK.�!	H���, ;�;�;���!�rˁW5��RE'�1��-pKIP_SKP���H�:"GM	_�ZERO�O�@E��`�����2�ǿ���2Nh�ˁ�5E���3��� @P�P�@��TDA�C�_LM��V��APRO�����#9DST��T�@��
b1K�KcF���m@	PʂEL�S��HjFLf`��Fgʢ ��y�F��J�I� ��`��d
[� US4�0�1V,\)TEX2]TX � ��^�t\SxZ�[�����6V��0X�� f��W	!�QS��1Q҃TD�aB����C`�B�	R���INj�CD����Hp����W0��yJhY RQ#൐0�Dek�Е�TUkg�j<u0SPE_WR@` �WEL�-�lY H�ICKNEzX�lTH29$TCPz�Uz?1_FCGA�x-z
�FGFL��$AUTCNT&�PAV�sJH+Bg��jq�����#CMPSSCA9 &�Cr0M@L�tu1FT��vS�p������@�C|DOTQ_�F�q�I�z���|�SMW��y�)��+RV����S�rh���) ��TP����C��EQ�1h����%0a����AF���𾍈FCTRLc�HI���GM,E1E��>bR#� ,AM���4D�SB^!�!l����#C�HVERACTI�V�#V�1��j�QZ ��#�!�!8��1w8�0��Q�+QQ�EQW8�FL�C^%8�3�A%0�Rh40U�GR�P�0.i�> x�C@LJO L�t!����	�
RE��LpdB����X�Ah�? �, $PGEA�PPL_F��d� �2=�Ȕv�> ���ҠSYSAT���i�@ `��!2�h3Vrh�ZpHRIZ�P�ET.�ERLM���E_DFL_���rI�DN����	�&`� TQ%��p��C}Dh�A @ ��v�UN٥EVELp�MA_�� HR-PU��s��qSEdq���F;  B	A�o�p� �1�qP���ER"VrLLOW&��DS_���Mb���SCRPL�����B&௸ƶ�Zp@� ��CH����1�"�����i0O \!�
��%�ݷ����Of�ROA_2G�=�(�1��9�M�M�������E��Q�v1SI3GNڢ��IZ,A@$�H��Y�P@�_�!x�C��*�$FO��DETAIۡ�r6�����HRONIZ���W2���qN/ _!PI �#��T!!b�?OAD_KA��8����y��i1"ß�FR8vP)�RC2Pn�dqzB��n_2��T0.�rSGL�A( `�@7�/@9�6�I �#W(�� Rn�REѡy��q@
E�u��n����A��VsXǒdC��l�p��tQMV2�U*�(����*ⱶV娲HO_P�s�P���q�
T|�A 8 Op{�I���q@������MO�I��P�r)�e �pSWI����Tp*�zBO�!SC�s��uN�@�p��!,�f�[�d ���0�LY��GD,�[�E�VNd����T0`L�MWR�ӌ� �$WT�q�v��Q�Pݣ�a��Jq'��u����GDIAG��X1�Ş��S'�I�`�RVI�I`p $DU?MMY166.%GDID���@&PHЭ�&N�cC�CD �p�0��4a�p���
h�<���NBPM�0�LM/q ��¿���
����VfЕ0߂Q�H�O��S��PEMP|�q��ELYWL��'DEF�f-�K���2�de�t��1��SDCL�iZsv� �P�2�TPZ3�!���TBL�঳HKY���UPW�POP��W[�v0% ED1>KNB_AR��>�ߠ���_��30��WpOPB_�$���/q��o�A��p�PD���ӍpH !� ��g,Х�? �S�q��)�KY78_2S���J� �[2	�_�AR7R_S��$�`�0�RS.��B_DB�q�2k�SGFI�LSC	q@OFF����TE[�� ����V�pPOm�F��C� r:9D3�:9FRO!�"�3?Ÿ�� R�s�5��uFCRQt�WT)MJ_�WېM�"��Nh`WT_~%�4ݳ���؀�U�FN_KaEY��S�N�AIP���WAVE|�P�W�L��*A��(CC!U,T"� /�N�#�2p�]HTP�p�ScB��p�_CAIRGAPS��FM����$��IS$��q�f�pDIH�CDO�H ���J��B��
U .�?��a !�p�sa��w�.V��DZ�C p� $UGA�PX_4GNcfQ�nU�A�G_��0��Gۣ�!�Vp�ЪT��O��[�D A��Q�u���_i�+�PTNOTRES�i5TRYd�-�?�a2- T��OL���F΀US�0��Tp�D��P.�`b�dXH ��fFL"�D-��|�FLA��TOU�AG�CKB���bEB�gM�p|��uB�|�Yp�AU_WI��T$6pcs���:Ch��#��Wb�DE��x}�c�rrSB_C��IM_PN�3�t��% ���qĢ�x�b�u���U��-�ERH�4SPT���tG��T~ �PT�e����VIC�P#R��ySP�QAV�Š�Q_���G�>�XBIAS4���p�sMPLd��d�`��{�h�������LNL���٣\0��`MG�P0{�ӈ�qS��0LMÆ�0���p����#����`! _��_�i�0CH&6�$���4&��H�"pU�MN��4PA��SW��Hr����0���aN61$�'��_�A@`�������W��I@OX��\�E�2G��~#d#��p$k�Q(aYuINC��AR�$9�v�tP�UP�WRHqG�?��0���c�Q�Vp0� ɠ�S$�0��Sא�TI(������JH�P)1����R<ذ�dDEBU5�;g�9�e� ��[�F� t$�1!�X�6��DY{CSK����8�va�IM��&�HCAS�>���"�RH&�o�BK�0F��0��`�������p��OBU���TM_s�!ⶳ�?RQDIFF"̴n��RSH۶ST0� P�ց^��!Է~�����������pKIEP��E�@1�=�_�p6�_D��)p�T�"�M��O(�O_ �2�9@OS���J�^��V_LE �Sq� F��[���T�D���d���Aq���TT�A��AVG��Ӱ�ĕ����
և����3�E��¿�ME\�f`�Wީs$�ֆ��q$���sK=Q��F�RT��~�_�P�`%���W��^�qrCND �፱qr��ڤ�������FL������מ�b`�D���s�SO_�<|B�1D4AC_��GNj��j窰_0�� �k�XЉꆰj�0�`k�Jտ��溂WT����w�LW�j��C�RR4AX��GN �%�����%�O��@�.�AG1Q�2%��2DX�p�O�PS��4�_�T���0����ЎSD���P�4�K�P��cTQ��N/�BK��xr����REDU�´� �q4�LW��P ǃ��qq��=��w`2ep4!p�LM�����m
EXP�p��A�BN@�c�bGVA�)`�P��� QCLB0��o���Q`$l`��p4`9N���OVR1��VG����q5`�B�9�EXEDN�TQL���V%UP4[���p��� �E�rU��Ú��<�}P� �SR"�>[RG x � ��@^��e����^�Wz�������PRG�_NP%�X�_1L��QQ�`RC��gH ��:�SPN!'ALIC�B��@y!� ���"���O����&������y!MTN��'LBD2 ���YZIՂr���#e�l5�PEE0YP�+�n�����INI����RSQ"pV�I� NT��0'p17�'PANEiPQԠ�o���P0�4X�@ I �¿����y�� �4�����28�T�0�5��T!�EQ:�^!IN�DEq�^)�F��V� <�HICK�NES^�<�XA��RV*ä�.����"p�1�94_p#p8��CG�HK`7��CG�Ѳ��OK2��QVT�`�#`��G��RB��17 ��JV!�P4cf`�>b
Dm
$�:@G� pT�_EQNO ��3�� 7�1��qX^a���� _v}F_LWĵqR�V�T�U�G� ����&\�!��T���cW� ��s�
Vn�P `r��6aqx��5K&:@�H�N2ap�#HOCGONF0��WB_�P2�ybAN^���Y@G�x�f\Fu�FLTRU���5D9pDO��P0\��u�UPU�0����k�bLW�k�h��RQ�c�b)xr�c"w <x�d��g^v�d^{|u\�p�MOD�#A�`@�nS��Tn�'PX�3$dW�p�rX�`S�TE`�TDCF~�J � $� ��g�}���q��{�u�&��OU(�0�W��v�IP� IZE�c_DH��l�PM���z�.�TD�� �RT)PG�l@Op�Z�����AT�PO���3"��Ԑ���s��K �JQe�ɑ$DUcRA�0䃿�DI�����9�ㄖ��j����9�ᆶ�ME3Q�$r�"���z�RE�V�Р��͂�L� 1�0吆�|���o�Z�o�j�U� Wf0}���I|���Q�L�<��|�ACTV�I�:�2ACHnB��0EXCf�$F�04{��6ːXIS:���1}�>��� �V�^�B96=����2����C�@�Н���T��FC栲���岩���ALE� ���W�FAUL���aI=�b���� LL. @�!3���E����2K� �����"��R���=�d v�}�Z�_C|�u@s��Ph&�ŕ�L AT�����DRO!�>!�u�݃���� G��ɒV��'��/�Ŭ� �\2HKb�M ��FL_E, I�	�`�P.�Z�E�Y�SW`� �v�� B������ȝ���DUMGMY0ƀ�"�0����Ǥ������0BII`��E����tG"��Dİ� ����IP�f1N 4 9@�1 �1A�PS. C ��C1��^�\2M� T ?O� $2ѿ �t�0�TE��ENS��Y�	���0������I�V��d��M_A����1���09�������ږ�F͐��O��Р� �MP��R�_AI��,�B5�AIF'�M6��u�9�<���_GIA��L1TRCPT��u�{�!_�p0�����S���ю��ALA�Ў��PM�. TAӴ�@@K�I�/�OV��OLCRx������ULST����2�4�-Pqԫ�?P  �y�o O[3RY-�f1Q L�p%� ћ�p�����-RLON��p�>WbA� PSH�!�Ȱ\1ZC�tR� � �@G0��uA�� ��%�������(���vAF�LSBK\��ȱZCD�L8�,���3$� F	���)��h`���䚐��B������PT�Q1�� �Hz@��TQPERASz@#��3� ��Fz� ��Ļ����0����DW���0��NLM_ZRO^��P�����7P;]�tZ}Cc4S � ��D�AU���uB�!G� ����LZ� 0�V> ��GN�2��ΐa@`�38J }$\1CAPITb�_ T ���M�;�pIAG�0��|��9$MEASC� H#9$�p$��PT�B��NBL�@A���!L܉R��NOM$�OL�1���'H��OL2�(2�%1$���$�-U����#BQ��$BU�Ff1U� $/WRTRA�YN$0 аC<#)/;/X%J(�1xN$T� WRFI]�X{6��|1MO��0`쀍5�2�7yARIŁ�M%��6�1�5{5z �ė3�5�5�:�:�4� ^ �4�6�4�5J!H�dfD��/�(Z��� ��qV� A9R�E1P]`�A��AUT�O[aÃdUMRY3FI�`��AK���GgWEAb!�2TU �2T�5#WY�6P5�`��UTUUk!1_�Bd�Cl 2yX$3A_:WAER�]N�!=�oK0FER��U�TD��V3�R}O�AD��-�'D�!M�0#W ���4;඗`/r/ �/�/�/�/�/�/�.)�A`4X �ۀ?'?0Voy�B���VG`u]s 9vhs9v�o�+��A`�qYX��ah�O�K�O0�K��/�B�Wgq��u_�_�_�_�_�_�VX��X���QX$LIFp�������WLDǄ��o(o�wSY��Z � 	$SG(�p��M>aA�d+��DINC�OO�YESCRN=�T�ޅ^�ޏ��+MWTC�W�[{  WELD<�_���NGLƲ��T�\��ә]����X�]3 <<Џ�URƳ��'PRA��2C{�C�wHEC������W�^ ��$䕉3'[ n�y�\}���F�p]��I�W�_\����y�^ ��$���Aΐ ���[���n�]n� ]�����SIONè�  1N��$FC�ONFI�G  ƥ�]P���GRP� 3�0 �	 �E��	 O�`�r�;�����Ŀ ���ӿ��k�B��f�9�uχ���S��� O��ω����<��� ̠)�z�M߉���߭� ��������A#�J�  ƥʢ��Ӡpgߔ�ߣ�I�[� ���������#��� t��k�>�`�`��f� ����������h���% I7m����� ��������! W��cwF� ��z�.//R/@/ v/d/�/�/�/�/�/ �/ /?(?�/`?�/�? ?D?�?�?�?t?O�? ,?&O�?\O�?�OnO�O �O�O�OO _�O"_�O .OF_l__�_�O�_4_ r_�_�_�_�?0ooZ_ To(o�o$o�o�o�o�o �oBojozoP&\o t�B��o�b� �(�� o^�4���� ����܏ʏ ��� 6������~�T����� ��p������4�� V�,�N���b�t���D� � �
�����.�d� v�Ư֯������п� ���J�<Ͼ���τ��Z�|��$FC_PDATA 30��] �  � 
Z���L�
����&�8� J�{�w�3�OФ�V�� �߷���g�����#� 5�G����ϐ�Cߴ�� ������� ���-�V� Q�c����������� ����]��
�<�\� ^p��ߺ��� ��J�0( ~��|�Z�j� //*/8b/t/F/@/ �/�/�/X/�/|/�/�/ &?8?L?��??d?\? �?�?�?�/O�?�?4O FOXOjOO�O,OnO�O �O�Oj?�O2_�O�Oj_ f_x_�O<_�_L_�_�_ �_o�_@o�_$ooto �o�o_�oVo�o�o (6o`�o��� ��V�z��$� 6��o����H����� Ə������܏2�D� V�􏎟��r�l��x�hø�FB 3��>���  �x� G�2�k�����v���ů X���*�����8�"� \��X�������P�ڿ Ŀ�Ϧ�4�"�X�� hώ�xϲ�H������� ߦ�0��T���Pߊ� x߮�H��߼����� ,��P���`��p�� @���������(���L�^��STAT �3!�] �Z���V������� ����	B-fQ �u������,6G� Ue�����) l������g/��/xv/�/�*�p���/ �/�/?+/)?O/P?�*���Z?]?�?�?�?D�?&(�?/�6�?�? �/?]O?9cO iL�4^�"�7���O�� �O�O__*_0_B_x_ f_�_�_�_�_�_�_�_ �_o>o,oboPg�~o �eZo�o�o�o�oLo�o (~�o�G	gw� �����	��� �-�c�Q���u����� Ϗ��ߏ�=�o�oM� �s�G����3ߟ ��ş���7�%�[�I� �m�������ٯǯ�� �!��E�3�U�W�i� ��m�+�}�翩�ѿ� /ω�S�͟y��cϭ� ���Ͽ�������)� +�=�s�aߗ߅߻ߩ� ��������9��ſ �A�C�k�{���#��� gϭ����G�5�k�Y� ��}����������� ��1UCegy �����_���- c���E%� ���/�)//9/ ;/M/�/q/�/�/�/�/ �/�/�/%??I?7?m? ;��?e?�?�?�?�?�W?O3O�?�����$SGATCS1� E]T�@�B
�@��@�@��G�O�K�O�O�DA �  @��B�D� T @�@BH�D�  CT#_5_�B�O�^_�O�_�_	R�@B�P  =��w�>L�P����@oE2xO�O�_ot_ *o�O�O__�o>_�o��oo�o�_�_�_CS3�_�_�o_�o�=o Ooaoso��o��r�7��o}CFG �1E7q�c���-�9q�������-�9s��-� (A������� �&���<q,�=�f� r���9q�����r��������  2����@�c���������0��f��sp<r`�qY�{� ����̅��܉P�ޏ(� ���¯8�7O@�C ���������̟ޟ� ����¿5�c�u�� }�ǯ��+�a�ׯ鯃� ����C�U�g�y��� ������b�տ�Ϗ� �g�A����wω�#� �Ͽ�R�������+� =�O�r�sߡ߳�-��� �{�i����?���K� ]�o���������P���<qoAD}���E�� -Y9u�����IAGo1 -}BEq ��Si{��������TWZR�CLB1������d m
/��Aq4"-�_��pe$bU�q�S��F�p,e/���u�W3?�U�R�,�/? 4�/0??T?;?x?�? q?�?��/�?�?O�? O=O$OaOHO�O�O~O �O�O�O�O�O_�O9_ K_2_o_�_�U��_ �_�_�_�_o�_,o>o Po#oto�oYo�o�o�o�!�__�o
�o @R%v�[m� ������<�N� !�r�����i���̏�� �����8�J��Z� ����Y_��ȟڟi��� ��4�F�X�+�|��� a���į֯�����߯ �B�T�'�x�����o� ��ҿ�������>� Pϟ�tφϘ�'ϼ��� �ϳ�����:�L�^� 1߂ߔ�g߸����߯�  ����"�H�Z�-�~� ��c�u���������  �o�D�V���f����� q���������
�� @Rd7��m� ����<N `3��i��� -�//&/�J/\/// �/�/�/w/�/�/�/�/ ?"?�/F?X?+?=?�? �?s?�?�?�?�?OO �?BOTOfO9O�O�O�J
�o�O�OkO}O_(_ �OL_^_p_C_�_�_y_ �_�_�_�_o$o�_Ho Zolo?o�o�ouo�o�o �o�o �oVh ����?��� ��.��R�d�7�I� �����Џ��Ǐ� *���N�`�r�E����� {�̟ޟ�ß�&�u J�\�n����������� گ쯿��"�4��X� j�=�z�������ֿ� ��Ϳ�0��T�f�x� KϜϮρ�������E� �,߻���b�t�Gߘ� �߼ߏ��������(� :��^�p�C���� ����������$�6�	� Z�l�?�Q�������� ������ 2Bh zM������ �.@dvI �������/ */<//`/r/���/�/ �/I/�/�/?�/&?8? ?\?n?�?S?�?�?�? �?�?�?�?"O4OOO jO|OOO�O�O�O�O�O �O�O_0_B_�/f_x_ __�_�_�_�_�_o �_,o>ooboto�oYo �o�o�o�o�o�o( :Jp�U�� ��� �O_$�6�H� �l�~�Q�����Ə�� ���Ϗ�2�D��h� z���_�������� 
�ݟ.�@��d�v��� [������������ *�<�N�!�r���W��� ��̿����տ�8� J��nπ�S�e϶��� ���������4�F�� j�|ߎ�ݯ����S�e� �����0�B�T�'�x� ��]���������� ��,�>�P�#�t���Y� ���������������:LU�$SGD�IAG2 ����s]% B�U�	�������"�TWZRCLKB1,7d@�+c
0O� AO   B�!b"�@���,�7J� ,� ��ր?�"� ,��5/��Y/@/}/�/@v/�/�/�/�/"
"/ ?�/7?I?0?m?T?�? x?�?�?�?�?�?O!O OEO,OiO{ObO�O�O �O�O�O�O_/_A_ _e_w_J_�_�_�_�_8�_�_jĐO)o ;o�_Koqo�oVo�o�o �o�o�o�o%7I mR���� ���!�3�E��i� {�N�����Ï�O��� ���/�A��e�w��� \�������ϟ���ڟ +�=��"�s���X��� ��ͯ����֯'�9� K��o���Џ����ɿ X������5�G�� k�}Ϗ�bϳ��Ϙ��� �����1�C��S�y� ��^߯��ߔߦ���	� ��-�?�Qu��� ������������� ;�M� �q�����h��� ��������7I m�d��� ��^�3EW� {�`����� /�/A/S/&/w/�/ \/n/�/�/�/�/?? �/=?O?"?s?�?�?j?�?�?�:
o�?O�? �?GOYO,O}O�O�OtO �O�O�O�O__�OC_ U_(_y_�_�_p_�_�_ �_�_	oo�_?oQo$o 6o�o�o �o�o�opo �o'M_2� �hz����� %��I�[�.������ v�Ǐُ�����!�� E�W��o{�����.�ß ՟矺����A�S� e�8�����n���ѯ� �������O�a�4� ������|�Ϳ߿��� �'�v�K�]������ ��x����������#� ��G�Y�k�>ߏߡ�t� �����߼�����/� U�g�:���p���� ��4�	��-���Q�c� 6�s�����~������� ��)��M_qD ��z���� %�I[m@�� �����z/!/3/ /W/i/</�/�/�/�/ �/�/�/�/?/??S? e?8?J?�?�?�?�?�? �?�?O+O�?OOaOsO ��O�O8OJO�O�O�O _'_9__]_o_B_�_ �_�_�_�_�_�_o#o 5ooYoko>o{o�o�o �o�o�o�o�o1�O Ugy���� ����-� ��c� u�H����������� Ə�)�;��_�q�D� ��������ݟ�>� %�7�Ɵ[�m��R��� ����ٯ���Я!�3� �C�i�{�N������� �����̿�/�A�� e�w�JϛϭϿ���� �τϖ�+�=��a�s� ��Xߩ߻ߎ������ ��'�9��]�o��T� ������������#��5���k�}����$�SGDIAG3 �������]V�B� ����������%�7S�TWZ_RCLB1>
]"hdq\�	
a�~� A   B� R�bS�@�� � ]T��h��,� �������?�S� ,��f�ϊ q�����//S�
SD/�h/z/a/ �/�/�/�/�/�/�/? ?@?R?9?v?]?�?�? �?�?�?P�OO*O�? NO`OrO=O�O�O{O�O��O�O�O_&_4Z��?Z_l_�O|_�_�_ �_�_�_�_�_ o2oo VohozoMo�o�o�o�o �o�o�o.Rd vI����� �?�*�<��`�r�E� ��������ޏ��Ï � &�8��\�n�A�S��� ����ڟ���џ"�4� �X�j�|�O������ ֯������0�B�� f�x�K���������� ��ɿ�,�>��b�t� GτϪϼϏ������� ��(�:��^�p߂�ѯ �߸�G����� ���$� 6�	��l�~�Q��� ��������� �2�D� �h�z�M��������� ������.@��d v������ �*<Lr� W�����/� &/8/J//n/�/S/�/@�/�/�/�/�/:
G_ 0?B?�/�/x?�?]?�? �?�?�?�?O�?,O>O PO#OtO�OYO�O�O�O �O�O_�O_:_L__ p_�_U_g_�_�_Q�_  oo�_6oHooXo~o �oco�o�o�o�o�o �o2DV)z�_ �����
��.� @�R�%�v����_���� Џ_�����<�N� !�r�����i���̟�� ܟ���8�J��/� ����e���ȯگ���� ��4�F�X���|��� �/�Ŀֿ������ �B�T�'�xϊϜ�o� ���ϥ�������>� P�#�`߆ߘ�k߼��� �߳���e�:�L�^� �߂��g�������  ������H�Z�-�~� ����u���������  ��DV)z�� q��#��
� @Rd7��m� ���//�(/N/ `/3/�/�/i/{/�/�/ �/??&?�/J?\?/? �?�?�?��?�?i?{? O"O�?FOXOjO=O�O �OsO�O�O�O�O__ �OB_T_f_9_�_�_o_ �_�_�_�_oo�_�_ Pobo�?�o�o�o9o�o �o�o�o(�oL^ 1C��y��� ��$��H�Z�l�?� ����u�Ə؏ꏽ��  �ooD�V�h������� ����ԟ柹�
��.� �R�d�7�t������ Я⯵�ǯ�*���N� `�r�E�����{�̿޿ �?��&ϵ�ǿ\�n� AϒϤ϶ω����Ͽ� �"�4��X�j�=ߎ� �߲߅����߻���� 0��T�f�9�K�������$SGDIA�GCFG ������]Y���� �����(��������G?UN1 5��&���]� BV:�D�� )���t�@�j��Z�?��  AL��A��&�B��@333���C�@Y�����#K@����(C��A�ff��2C���A녇�9C̿�A4�͇�?�C�"�AK��?�D�Af��?p��2&�!3E�ad���
>܃�@?�`��<g� ?����� ��R�����:E�ᱱT��O�,���V�Apτ�ss��?�tv
,��L����^�?E��� ��cT  _��p/�/�(7�/@[�_�#��"��>A$/?�2���A����
Ph%�/B?��0?�m?�]"
Fo�rceCheck��p��D"@���2(���r d��d�9\��3 BHf�1[�sD]��� �1�<�B�� 1�2�s�1�11DB`-O?OQOcFn�t"
 �I�O�O�O�O  __�O6_H_Z_l_~_� ^�d�14
�T	���D��YA2�0P#�_�_�T�Z�q��72o  8�5eh8"  D����MG=����B�D��_>�� >���$eHo�h�,@t +�9>1:  ��h��	r �4��7�om�h�� hc��D����%T�t!\D�+�����1�C���?�?ff���s�5�Bu�40�& G̖��_�S�w��; ��r�J�# @��C�r  F���6�Q��P�C hqL"ip�1?��>`  <,T{J��� �W�: �j�F#��R�!��07-JU�L-21 04:12�\�i �/ď֏@9���u!��1�10���~�?�p�B����6�陚A33A#��R�d�v���_J���沟ğ֟
 ������!���E�W� i�4�����r�ïկ� ����/��S�e�w� B�������ѿ����� �+�=��a�sυ�P� �ϻώ��������� 9�K��o߁ߓ�^߷� �ߜ߮��������G� Y�,�}���l�����@�����R�22�〔�)5t��^J�!Z� �t��BlR�":�$��o����48!?�0t$�!F���@�1I
J@7fff(d=�pD%� G �D�
@
���T(�T+!_a+!2��=��T���k�q�q'WF�#��i��(�!B���6�4�q�q��!��o$@�`�1�z���@y���$,�S���P�/P�pPF�N�q��h eo�P�1|u |�� c���S���34�rq� @#� `r�DH&�I-�1�q�2t/��/��rM� �*�/6�	��(�_��I�qq��'3I�$< �p@9H�*��UKKU0 ���a�1D�r��T1$�=�2)�2 � �1)T10q�=T?^�����A�#
?2r�3>  ��2I�$D�/���q1s$D������� X  �p cq1���!�@�Q?�O�@�N�a��O8�F���=8�-'_ _��d_v_��[_�_�_�As P�� ~t�Q����2�
6�084��1�Qe�(�J4a{�{2 / ?20f?�����o+o=e?�?��c<�Pb���pԒp]n���:h��M?�-Y�@��1BF��Zo�4n�I�?�0�|D��b6ffBJ���oF4:hȭ��?�0lH��bY�g�B�o4aBL:h�L�?�;L�>�a33B1F�=~F42�R,�>{:a �s>c`?�����  ��DC�S�S��P��� ������������Ǐ� ����L�3�p�W���Ȧ�Q�#S�*2ʜ�$�SGGUN2 �5�����]�IS��%C����QB@��e��B=x��AKprM� �DC�`�N�#K�E2C���L���L����L��"�HUD�甦f��*�唦;T��L^��D] R��n��w%P���hbʟ`�R3�.�>�<#S L�X�>�L�n���6^B�и�7����A�F!,#6_P�L��#U�#Y33#_�Ll��@zϊF��j�K[�S�lD+�5 c��� �� ���5�A�ۿQ��	�� +ʀB� ,i�R���P%���ߒT����'�<��
SUe5�	�P(�d`���SG�� ��S�3(��"���;� t��Qc�3P%t�������	��R��B
 D�\�n������� ��X�������"����d�A�s2�t	��������B���� @�T�0B�SD����,M��&����� (���?æf���� �S0 ��A�׵!Q$�T;� ���NR�S +@U���:0�!A6�<`W!�2!��?A�R{A{#��/��/�/�Q��&��*,�/�ߩ� ӿh?z?�_�?�?�?�?��?�?
OO/?��!9/`OrO���?�O �O�O�O�O�O_�O1_ C__g_y_�_V_�_�_ �_�_�_	oo�_?oQo $ouo�o�odo�o�o�o �o)�oM_2 o��r���� �%�7��[�m�@�R� �����������Џ!� 3�E��i�{���`���ß�,2��<�/�,�2m�/�Z ����F��j�D	3��?e��/�Fb��@e���
��@fwffA-=̮ ����������
@
	�l(lk!k!2,��j{�8��9�w���F�*�m{�/�B�$M�L�W1W1Ș�ؐ��ȡ@`��z���@y����`�~��  	�@q Y �~��}!b��	��a�M� ��  �]��P�b�a�;��P��״�"0 �$0 ������9���1���M�}!2�t�:�8�P"���!�d�ژ�!#�Ln$�#��c���� ȡ<ɠ���/�*o� �������������(� ��"1���ȱ\�(�Ͱt���}�Ͱ�������ߊA19��
?���� NA��Z3H��oߞ���!��� �!W2��/c���d�߆{�������ߡ 8/Z�����k!��`����Pba�A� P� "$�)� /�`�8�/�*{�֠���� ��0/AS ew������ �//+/=/O/a/s/@�/�/��)��/ݣ�B� �/,?[�P?7?t?�?m? �?�?�?�?�?�?O�?�:OLOg������nL��$SGGUN3 �5P�P�]�/�����C�@�v:B@�B��СB�nF�����O__ *_<_N_`_r_�_�_60ץ/��_�Z<���- �_�_�_oDo��#�th`�o�[�S�Q�V,����ۥ��o����ס0ץ�������l �V6�_����+�L� c�p��4oVo�� �xo�g�7A�j$� д�N0��_: %a��� 6x���w�r�o�������������Dd�l�� T��Y'�g� ר�Drt�0��n�� sע���w������Iw�(�
 �I  ��$�6�H�Z���~�@������Ư�OF~dT� 0��E�4O=�,Oa�s��Y�s ������Կ�7�2u�Z��йt�E�R��M7@� �����?�fft艬��0 $���ߧY���6; ��`����� @���bB��S�#�6� ����L��'�?�����d߳/�qߚ�7�pb���sе��K��kwo� �5B�T�f�9���p�����ߩ������Q��p�E�W�i� <�������|������� /��SewJ ������� +=as�X� ����/�/9/ K//[/�/�/f/�/�/ �/�/�/?�/�/G?Y? $?6?�?�?t?�?�?�? �?OO1OOUOgO��в2FC�a�е���|���Z �б ��Y��OQ�_���Ӂp�?	��t�FP@�	��S
�Q@fffAѳ=�RЍtfp�M��rp
@��B�(�sq��sq2�B��_��HR�S[��U�Fx��@���c�4��������<�4�Nk�lQ@`2üz��/@y��x�S"a?�  	�w���P�a"a�l!�P�b �a�cPd��j�p�nW �R�o|S�U#5{{d,ҹ� ���Zq2 �o�hݔ�v�a�}d�!с2���U�D No/��~HQ���Ԃ��p�Qo���lQ< mP���ߊ���T�S�� dbea=a=ae`̂a�DҀ�d��la �̂q`� >`!�q`��x�0���.ĸ��ݑE�
?z�D��P ��z���l��B@�E�y�l�[��� ��c���R(��L�*���C�1�;��Q���� \�y��?O����5O������oAe� EP����7���8��ӕʀ8�߆�{|���wq����y��� Կ����ӿ���	�� -�?�Q�c�uχϙϫ� ����������)�;�%�͓�߁S��[��� �O�����*��N�`� 3���}���������k��r���$S�GNRMCFG �36����]"���Js�O��ۢ�{U����|rۢ% ���ڤ����ȕ�E�rB�UT��yqk�>͐� �`�5`���S$�EXE� ;1�]%]�Vh��B� T�f�x�����������,<� �1������,		|��� x/(/:/�^/p/�/ /�/�/�/P/�/ ??pQ??Q �Q L?�?�?�?p?�?�?�? �?O�?5OGOYO$O}O lO�O�O�O�O�O�O_ �O1_ _U_g_y_D_�_ �_�_�_�_�_	oo-o �_Qocouo@o�o�o�o �o�o�o)�oM<q�V{�r>?�c��0,��� �%��I�[�>���� t�����ُ�Ώ�!� �E�(�i�{�^������ß�PFB1 <1�������?�ҟ�2�O�+�������ƯY�3h���ί���A�ԮRSF1  �A6������� ¿Կ���
��.�@ϸR�d�V�1B4i�p{�����u�SF2i� ����0�B�T�f�x߀�ߜ߮���������2@�Ϝ�-�?���d�3�� ������������
��.�@�R�d�V�3@
�����s�d�Ih����������� ����*JN` &u���h�������A`�MSG��2�FXdp ��W��/�W�CFG @" 7T -�m%r(��q�r  (�t#�q�$�!/%b/t/�/ �/�/�/�/�/�/3���XDATA ?�����_�/ (^ $1�?��8 ���2�Ϥ1 W �S�0'�3�1�0<�<�0�V�H��?�³�c!��0�1�������)2�a�m?�  E�M�@�o�lDc���p1�5<���?�!���8��!@A5�R�5�Xv7�� C�S�\DDb��aA�1����`TA�<�?�?�?a�O�!O3O\EDa�KF��ff�A�?�O�\O bq�;�.��@@ 0Q3-P�﻽.3AP�����0Q��1'Ĉ?S3D?%��p#_�5_G_YT Y�7����캷��j0ʺ7�; �"e� 2Ǻ���kj0�EZy��E�� đ�� \Y�_�_�]�2`�1r�7�,b	[ D`�!gKo]mEmEo�i!<�b	PD�  �aQC   �a_�d�l0�v�o�o�r�64�1��1�hq��aaeE~ĕ�r�prpi@�	m@ $���?�{�L��Ӂ<0�1 |v\�!J���y�vW^t�1w/ ,8j (|�2�^|�?B|  <P��mA]dPh� q� A Ad�v��	��<�� }A����4n�	 ��̂p�
�	.�  8�=�?�;@U@t�d�Z@U��?����4mI��I�"���7\q�T�/��\�D���oP����R�<o  ��H�Z�l�~�0����=�̩��_dQx� ����� �"�P��� >�`���8����n�� �,ϒ��^�ȿfϔ� ��Kϩ��ρ����� M�7�A�s߅ߗߩ�K� ���������#�+| Z�l�^��*߬�/ߤ� ������wТa��X� cz�i�it��������� 4�̀c�	��-��Q c��|���r�� ̟V�l��2> x�����ȯگ /�� �:/��B/p/b �/"/�/�/X/�/ ?�/ �/:?L?�/?~?�/v? �?�?l?�?�?�?�?2O O"X?bO�O�O�O�O lO~O�O_ _2_D_:� L�~_�_R�d?.OPO�_ (O�_o9o$�6�H��o l��o���o���o�o�� #3YX_}`�O ����$��1� �.\�j�t������� ȏڏ��	����_
o ,of�on�����ğN� ��������,���T�f� x�ޟ<����¯�Ư ����(�ί0�^���O ������ҿ������ (�:�L�^�p�f_x_�� �Ϯ_�z������� D�>oPoboto�ߘo�o �o���o� �O�: s��ϩ"����� ��.�P�9�$�]� ��� ��������������� #f� ���V߀3 x��bh��" �*X����
 h�@�/� /"/ T/�\/�/h����/�� �/�/?"?�/B?T?f? x?�?��.?�?��z 8/�/(On/ O^ODOj� |ߎߠ��O����__ �?:_�/j�{_f�_�O �_�_�ON_ oo$oZ_ ,�eoP��oLo:o���_ �o�o�o �j�3�gy�tg^W��lr���2�23O�sO�KO����r�   ��� �J���R����k�*   �����$�r����l� 
�8�2/,�n�P�&������\Z:��[��0�@n	�P�?��7�Q��al��LC�@��Џ������I ������1�ud̢�?�?S�: F���?\�ʟL�ϟD��f����O�o�4 =x�O~o(�B|  ��M@�/0�]0�����`���@b�^x�@n>���P��)�φ_»!K����ԯ��0�o2��éo��<�,���?��`�@m972�xTo��xe�QGO�Q�Y��ހ������ �������#�5�G�Y��@�����v������ � ,,		 �ᴥ ����.���_� 5�����������[� ��������?��� M�%����!�� �=�[�Qs�� �������/� 	/7/]�E///�/ �/�/��/�/-?G I?k/�/{?�/�?�?�? i?�?�?�?O/O�?g/ =OwOOoO�O�O�//? 	?�O%_??A_�?�Os_ �Ok_�_�_a_�_�_�_ �_'oo_O%oooIoo �o�o�O_�o_7_ U_[_�ok�o�o�� Y�����1�Wo �?�y�������o ��/MS��Ï u���}��������ß ����)�O�ٟ7�q�� y���E�ߏ����'� E�;�]���m���u��� ɯ[���뿑��!�G� ѿ/�i��aϟυ�ׯ �������1�3�Uϳ� eߋ�]ߛ߁�S߱���������:�Q��$S�GSYSATUN� @(�]�;�w�		�o�T�CD Ab�z����z�S�CFG QBb�S�t���c��i�������y��R���D����x�xv��� ����%�r�v��E����G�=���4 4�Jء����� ���>R� �@���]�"������2�����?�y�
y� 
��	�u�d��,�#�F�y�%�����0S�S�4����`����C6:\E�VENT_SPO?TWELD\��@
.@Rr���P��%�I�T�D��C��������TCH !D��%����/�����r�%��U����m/������/�-�������@�v-_"C��/�&�W:��E�  bw��� L)25( $�Z5������EXE I(�]%��?�?��?z/�?�y�ZO ��-DJA ?KTN q?xO�O�O�OM�O�Oo�,�_,_>_P_$b_s]�?�WgO�_ �_�_�_�_o??NCo�'H��wo�o�gao �o�o�o�o�o#�o GYk9���� �����1�C�� g�y���Y�����ӏ�� ��	���?�Q�c��  �ϊ��ϖ������Ο ���>�(�b�L�^� �����������ܯ� �"�h�
�_t���b������$ ��f����Uf�y4 u���?ֿ���>)� `o2�D�V�0�zόϞ� l������ϴ�
��.�@��R�d�v�ƿ�7B)j�p �����@1?��@����� (�|�&�,�2�4�F�� j������t�"�� �(�B�L�^�p�>��� ���������� ��$ 6H���r��~� ������&���2DCF�J������ ����&
g4g4lC?�4DS�2K"; ������!L%���\I���9/ K/	/O/a/s/!/�/C�SET 2L"9i0�l>5? ?����FNH@@>6598<>;=>L��x8>�EHK� 1 M�-Y��$�% � @#x�@��:@��A"���>?OF�0?���?m��?�?(�?��OLO�H�F������VOS<`�>Ͼ�����TAQ4�72�<aKyO�O �O�O_/__?e_pW�O�53�O�Op_�_�_ �_oo�_T_Pox_�Z�IPCMP N��@M�aSO1 P�]{:C�����A  =�9=X�a>,1�a�1@md�=���i�i2�o��o^�o�o)~3 ;M�q����(�OFFEXE  ��;�_ARYO�UT Q�+� D�*���:@EUN�F1  �; �By�nD��Cz  ��p���Bށ��^�DvpC��E?W�A���1Ư�B4��ˏݏ�E�.��2�l�x�t�P� �e�ş����3���� �ڟ쒢��a�%����I���;�#R�!�  ��^0�� @e
 �  D�^w^[r���>� ���ѥ���ɯ~�T�� .�n���6���K���Ϳ ߿��𐪿�*�<���=��Gωϛ�+�MSAG��Q�������""��H�Q�4� �ϻ��#߃�G߻�K@f� T�0�%>��e�1(�أ1�1�1 �����������!�3�XE�W��&ZCKR�}
pd B���Q0�T�!Zp�)� ]���	�a 2�� �j��5!���W�S�^ �=�^88�|2���DTCAP�0	V�+@a|������a5 �!@d�c ����$�h�121-0�7-28 01:33:2�H=:? �{������DK�:E�! �����2�����[m:���|��� �I�)�!T�%�a���`���/1 ���",/�bnanaK,�<  (25:04QU�/??�� �@���1��&n?�?�? �?k?�?�?�?�?�/"O 4O�?OjO|OCOUO�O �O�O�O�O__�O�O T_f_��� �_�/�_ �_L+_�_�_o�_�_@o�_jo!o�o��3:? L?&_�o�o�o< N`'B_��o� ����&�8��� J�����Y�k�ȏڏz_ ��j�o$�|o2o��� ~�5�G�Y�k�؟����.��MTR��Y�o���� 2345678901C�k����� r��#C�U��������� ����y������^� ��$��90"� 4�����ؿ4���ǿ � 2�ү����Z�l�~� ��������`������ �O߫�,�>ߗߩ�I� u���e������	�J���Ͻ�SYS Z�	ݶ%�`�'��_MW�TGUN1 _�	��a �  \�������� ���>�P�b�t���� /�������������( :L^p��� ��� $6H Z�~����m ��/ /2/D/�j��2���/�/�/�/�/ ��/??1?C?U?�/ y?�?�?�?�?h?�?�? 	OO-O�?�?cOuO�O �O@ORO�O�O�O__ �O'_M___q_�_*_�_��_�_�_�_oT/��3 l/~/Ooaoso�o�o�_ �o�o�o�o�o9 K]o�(��� ����#�5�G�Y�  ��������ŏ׏n� ���1�C��S�y� ��������ә