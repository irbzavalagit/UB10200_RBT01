��   ��A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ������IA_EL�EM_T   �D$USE � $LINK�_NOD HTY}PC$SHA\�IZ]DATA �  �4�/HAND7 �< $3 3� � SLDIST�D $COMME�N� $DUMWMY3D �4��� �$$CLAS�S  �������"��"� VE�RSION��  1N��$� 3��"� 
  0��c��4  C��1r Ug�����/
��
/ � '�V/ 9/K/]/o/�/�/�/�/ �/�//#/5/?d?G? Y?k?}?�?�?�?�?�? �??1?OOrOUO�O yO�O�O�O�O_�O&_ -O?O_#__c_�_�_ �_�_�_�_�_�_4o;_ M_o1ooqo�o�o�o �o�o�o�oBIo[o -�!���� ����P�Wi;� ��/���Ώ��ÏՏ� (���S�^�w�I��� =���ܟ��џ���6� �+�a�s���W����� ���ͯ���D�'�p9�o���	NUM� V�    
