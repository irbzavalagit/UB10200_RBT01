��   8��A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ����DCSS_I�OC_T   �P $OPER�ATION  $L_TYPB7IDXBR1H[ �S2]2R4�$�$CLASS  �������Pz��P� VERS?��  �1N�$' 3 ��P @� �����
(�� ��� �������" �������
�����b� v�������j(���� ���� �*����~ �b�v�{/a	�/�"�~��!.���^/�'�/  �s61� uR1��sn1�s�1��s�1�s�1��s�1�2 u�1��sA�_?  A_���!��$"jE� �$�E�!!�(��E�"�$Z�E�#�$~��E�!$�$v�E�%�$� Q%_7_I_[_m__�_ �_�_�_�_�_�_o!o 3oEoWoio{o�o�o�o@�o�o�o��R1"�o���m�/Y ;Or61:O,s61VI� Jq61��fq61F��_C_CCL ?���  	�All para�m��
Base��Pos./�Speed ch�eck(�Safe� I/O con/nect�}R��`� �2�D�V�SIi��@{�ExtEs�top��ǀt�yFnceClo�sed��Rob�otDrives����AuxPowser9��T1-���KeySwitc�hU�2`���3�D�isabl#� Reserv��𞟰���sblM�ontSpaceI1���2����3����4,���5D���6$\���7t���8����	9��0���oׯ鯀���ǁ����*��	�Zero����ƁS_ignLaj�_�f�ch��~�x�����q�IO%�Tool�1SelԀĘ̳2$ӿͲ3�Ͳ4�ͲI5�Ͳ63�Ͳ7K� �oρϓϪϷ����� �����#�:�G�Y�k� �ߏߡ߳��������� ��1�C�Z�g�y�� �������݇O�{�m.�ES�PB���Always O3ff�.�FF̗F���Auto���T�������D?eadman�ǁtyBypas"�� CellP�rimǁʙ' Zon����+�C� [�s����� ��N�ԥ������*�?����C��j�d{�L������m�edõ̿޿� ��&�?/J�\�% �/�/�/�/�/�/?? @?;?M?_?�?�?�?�? �?�?�?�?OO%O7O `O[OmOO�O�O�O�Oh�O�O��N�  ��	_��;_M___q_�_ �_�_�_�_�_�_oo %o7oIo[omoo�o�o �o�o�o�o�o!3 EWi{����`������SIh� ��#��f�x������� ��ҏ�����,�>� P�b�t���������Ο �����(�:�L�^� p���������ʯܯ�  ��$�6�H�Z�l�~� ������ƿؿ����  �2�D�V�h�zόϞ� ����������
��.� @�R�d�v߈ߚ߬߾߀��������*�5�P�%_�W���24V>��SFDI���� D��\��t���� ��� _/�A�j�e� w��������������� B=Oa�� ������ '9b]o��� �����/:/5/ G/Y/�/}/�/�/�/�/ �/�/???1?Z?U? g?y?�?�?�?�?�?�? �?	O2O-O?OQOzOuO �O�O�O�O�O�O
__ _)_R_M___q_�_�_ �_�_�_�_�_o*o%o 7oIoromoo�o�o�o �o�o�o!JE Wi������ ��"��/�A�j�e� w���������я���� ��B�=�O�a����� ����ҟ͟ߟ���'�9�b�V�Od�v��O�ﯣ�ﯣ�ﯣ�� ���ﯣ���&�`�Q� c���������ԿϿ� ���)�;�d�_�q� �ϬϧϹ�������� �<�7�I�[߄�ߑ� ������������!� 3�\�W�i�{���� ���������4�/�A� S�|�w����������� ��+TOa s������� ,'9Kto� �����/�/ #/L/G/Y/k/�/�/�/ �/�/�/�/�/$??1? C?l?g?y?�?�?�?�? �?�?�?	OODO?OQO cO�O�O�O�O�O�O�O �O__)_;_d___q_ �_�_�_�_�_�_�_o�o<o7oIo[o�ox�S�I����SVO�FFnoFENC�E�oEXEMG��oSVDISC��nNTED�o�OP�oqAUT=OT1L\r���<�MC~rC�SBP�
PO�SSPD_ENB�sjCONF_O�K�~F_IPARG_CRz�g����~��o�q_�o;��o=�y'�C_"�r_`��y 