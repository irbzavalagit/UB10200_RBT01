��   �=�A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ����EIP_CF�G_T   �� $VENDO�R  $DE�VTYPE>PR�DCODIREV�ISION>FA�ST_UDP �5 KEEP_IO�_AnSCNpO�PT` Sp $L�OADED� �C�C� IG�ED_wMOD�NET��EXPLCIT_�MS�$HIG�H_SPEE��$EN8qDS+CP� Hp �� �SPARE�4�&ONN. |� $HOS� �!B SC9ENA�BL$STA�TN _SZ�S�^TOAPI�OETrIgA�R]�V�BW&Mo�SC.�  7�CXQ�[�XX_���X_��[ kRs)%'wFLA�MUL�sTR�� C_O�6["TOD&ICi ��AS�Z 'EC�{#�#TIMVCN�� Z�&PAT � @$IDA_FORMA��!�&8� �"9"FIG^�"�2�+�!�$AN�ALOGI�  � 4OU� 8F�M�$Q�(4��$$CLASS  ���e1���.��.Z0VER�_c7  1N�$'0 �8�. d���� ���0�?��0���7/ ��4( �3�;@ p!172.19.A���?�4<���s;@> �1d!�  ectionA�BO�6�1 _L�:!�H12HO|ASS�W1 WTC n��OQN�DRI�G�J3��O|AWater Sav ?OQN�1�1�O|A(__TD� Dump on	4q_���OuO�C�_�SCapChan�ger1 ;�1 $�ka/_�_�J�l1Co�LReser?ved n6Qo�o�o�W@oRoApp/2-1 <@7�o�oP�o'�m2�a81�as��m3�a9@������m4�aA�A�S��w�Zol`�B����Ïf���k3�cC�!�3�֏W���JrDa�����F�ǟ���rEџ����7���*�FA�q���&�����l`G���󯖯��k4�cH!�Q�c����*�JrI����ӿv���*��rJ�1�C��g�*�*�Kqϡϳ�V�����l`L���#���G�
�k5�cMQ߁ߓ�6� ��Z�Jr0���ߖߨ�)�\ۺrO1�a�s����Z�*�P����������l`Q�A�S���w��k6�cR������ f�����Jra0#����Y���rTa��F���*�U��7�l`VAq��&��k1-5�aW ����/�ooK/ ]/ /�/$/��o�/�/ p/�/�/�O+?=?�/ a?Dfe�?�?�?T?�?�5�?OO�?BO�? �`:/{O�O0O�OTO�a �/�O�O�O!_�O�a? [_m__�_t?�?�_�_ |_�_o��?;oMo�_ qoo�jO�o�o`o�o �o��O-�oQ�o �J_��@��_�_ �	���?�2�*ok� }� ���D�6��oۏ� �����6�
K�]� � ��$�6�z��͟p�� ��'�9�ܟ�o�b� Z�����P�ѯt�f�ʏ ����A��f�:�{� ��0���T�fѪ���� ��!���W�i��� ��������π�ߤ� ����;�M���q�ߖ� j��߽�`��߄ߖ�ڿ �-���Q�4�Fχ���<�N��� !Spare�������1� ����g�y��.���R�����������$EI�P_SC 3����.� @�����  K�������@]�H����}���� �,>Pbt �������/�/(/:/L/^/�� Af/i/�/�/d������/Ij�+	�{4�" ?$�,�,|�A? S?���?�?�?�?�? �?�?OO+O=OOOaO sO�O�O�O�O�O�O�O@_�/'__K_�-����+9Rh_J�/?�s+uR)0,e/? �_�_e5>Q>_�?4oFo Xojo|o�o�o�o�o�o �o�o0BTf x��3_������rQrP0*��_�_n�_4+qP*0'2�f�_~���c7��
 o$oՏ�����/� A�S�e�w��������� џ�����+�=�� a�P��������.�@� R�d��'���uR�!�� 6�x���������ҿ� ����,�>�P�b�t� �ϘϪϼ�����w�� ��(�:�L�?ѯ�u �߸���]?��a��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z�ߞ������� ����k�}ߏ�@Rd ��=�߬���� *<N`r� ������// ����'/9/n/�/�/ );�/�/?�� 1?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�OW/�O �O__,_�/�/�/�/ �_�_�_?�_A?�_o o(o:oLo^opo�o�o �o�o�o�o�o $ 6HZ�O~m�� ��K_]_o_ �2�D� �_��_������ԏ ���
��.�@�R�d� v���������П��� ����N�`�r�� �	��̯ޯ�c�u� �8�J�\�n������� ��ȿڿ����"�4� F�X�j�|ώϠ�7��� �������������� f�xߊ�����!����� ����,�>�P�b�t� ������������ �(�:���^�M����� ����+�=�O� $ ������l~��� ���� 2D Vhz����� k�}���./@/R/�� �������/�/�/CU �/?*?<?N?`?r?�? �?�?�?�?�?�?OO &O8OJO\OnO�O/�O �O�O�O�O_/q/�/�/ F_X_j_�/�_?�_�_ �_�_�_oo0oBoTo foxo�o�o�o�o�o�o �o�O>-bt ��__/_��� w_��_L�^�p����� ����ʏ܏� ��$� 6�H�Z�l�~������� K]ǟٟ� �2�� ���������#�5� ѯ��
��.�@�R�d� v���������п��� ��*�<�N�`����� sϨϺ���?�Q�c�u� &�8�J߽�n�ᯒߤ� �����������"�4� F�X�j�|������ ���������B�T� f�x������������ W߽�{�,>Pbt ������� (:L^p�� +�=���� //�� ������l/~/�/ �/�/�/�/? ?2?D? V?h?z?�?�?�?�?�? �?�?
OO.O@O�dO SO�O�O�O/1/C/U/ __*_�/N_�/r_�_ �_�_�_�_�_�_oo &o8oJo\ono�o�o�o �o�o�oqO�o�o"4 FX�O�O�O��� 7_�[_��0�B�T� f�x���������ҏ� ����,�>�P�b�t� ����Ο���e w��L�^�p��� ����ʯܯ� ��$� 6�H�Z�l�~������� ƿؿ���� Ϸ�D� 3�h�zό����#�5� ����
�}�.ߡ�R�d� v߈ߚ߬߾������� ��*�<�N�`�r�� ����Q������� &�8��Ͻ��π����� �}�;�����"4 FXj|���� ���0BT ����gy���E� W�i�{�,/>/P/���� q/�/�/�/�/�/�/? ?(?:?L?^?p?�?�? �?�?�?�?�? O�$O OHOZOlO��// �O�O�O]/_�/2_D_ V_h_z_�_�_�_�_�_ �_�_
oo.o@oRodo vo�o�o1O�o�o�o�o �O�O�O`r� �O]_����� &�8�J�\�n������� ��ȏڏ����"�4� �o�oG�Y�������% 7I[��0��� Q�x���������ү� ����,�>�P�b�t� ��������ο�w�� �(�:�LϿ�џ��� �ϸ���=���a��$� 6�H�Z�l�~ߐߢߴ� ��������� �2�D� V�h�z�Ϟ������ ����k�}Ϗ�@�R�d� ��=��Ϭ��������� *<N`r� ������ ���'9n��� �)�;���/���� 1/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?W�? �?OO,O���� �O�O�O/�OA/�O_ _(_:_L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHoZo�?~omo�o�o �o�oKO]OoO 2D �O�O����� ��
��.�@�R�d� v���������Џ�� �o�o��N�`�r��o �o	̟ޟ�cu �8�J�\�n������� ��ȯگ����"�4� F�X�j�|�����7�Ŀ ������������� f�xϊ�����!����� ����,�>�P�b�t� �ߘߪ߼�������� �(�:�ѿ^�M��� ���+�=�O� ��$� �����l�~������� �������� 2D Vhz����� k�}���.@R�� ��������C�U� �/*/</N/`/r/�/ �/�/�/�/�/�/?? &?8?J?\?n?�?�? �?�?�?�?_q�� FOXOjO��O/�O�O �O�O�O__0_B_T_ f_x_�_�_�_�_�_�_ �_oo�?>o-oboto �o�oOO/O�o�o wO�o�OL^p�� ����� ��$� 6�H�Z�l�~������� Ko]oǏُ� �2��o �o�o�o������#5 џ��
��.�@�R�d� v���������Я��� ��*�<�N�`����� s�����̿?�Q�c�u� &�8�JϽ�n�្Ϥ� �����������"�4� F�X�j�|ߎߠ߲��� �����ߑ���B�T� f�x����������� WϽ�{�,�>�P�b�t� �������������� (:L^p�� +�=��� �� ����l~��� ����/ /2/D/ V/h/z/�/�/�/�/�/ �/�/
??.?@?�d? S?�?�?�?1CU OO*O�NO�rO�O �O�O�O�O�O�O__ &_8_J_\_n_�_�_�_ �_�_�_q?�_�_"o4o FoXo�?�?�?�o�o�o 7O�o[O0BT fx������ ���,�>�P�b�t� oo����Ώ���eo wo�o�oL�^�p��o�o ����ʟܟ� ��$� 6�H�Z�l�~������� Ưد���� ���D� 3�h�z������#�5� ���
�}�.ϡ�R�d� vψϚϬϾ������� ��*�<�N�`�r߄� �ߨߺ�Q������� &�8﫿��Ͽ���� �}�;������"�4� F�X�j�|��������� ������0BT ����gy���E� W�i�{�,>P���� q������/ /(/:/L/^/p/�/�/ �/�/�/�/�/ ?�$? ?H?Z?l?�� �?�?�?]O�2ODO VOhOzO�O�O�O�O�O �O�O
__._@_R_d_ v_�_�_1?�_�_�_�_ oo�?�?�?`oro�o �?]oO�o�o�o &8J\n��� ������"�4� �_�_G�Y�������%o 7oIo[o��0��o�o Q�x���������ҟ� ����,�>�P�b�t� ��������ί�w�� �(�:�L���я��� ����ʿ=��a��$� 6�H�Z�l�~ϐϢϴ� ��������� �2�D� V�h�z���ߍ����� ����k�}���@�R�d� ׿=������������ ��*�<�N�`�r��� ������������ �߽�'9n��� �)�;������ 1Xj|���� ���//0/B/T/ f/x/�/�/�/�/W�/ �/??,?���� �?�?�?�?A�?O O(O:OLO^OpO�O�O �O�O�O�O�O __$_ 6_H_Z_�/~_m_�_�_ �_�_K?]?o? o2oDo �?o�?�o�o�o�o�o �o�o
.@Rd v������� �_�_��N�`�r��_ �_	oȍޏ��couo �8�J�\�n������� ��ȟڟ����"�4� F�X�j�|�����7�į ������������� f�x�������!�ҿ� ����,�>�P�b�t� �ϘϪϼ�������� �(�:�ѯ^�M߂ߔ� �߸�+�=�O� ��$� ���߻�l�~���� ��������� �2�D� V�h�z����������� k�}�����.@R�� �����߬��C�U� �*<N`r� ������// &/8/J/\/n/�/�/ �/�/�/�/_q�� F?X?j?��?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__�/>_-_b_t_ �_�_??/?�_�_o w?�_�?Lo^opo�o�o �o�o�o�o�o $ 6HZl~��� K_]_��� �