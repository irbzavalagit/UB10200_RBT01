��  Ij�A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ����SBR_T �  | 	$S�VMTR_ID � $ROBO�T9$GRP�_NUM<AXIaSQ6K 6NFF�3 _PARAM�F	$�  �,$MD SPD�_LIT4&2�*  � ���4�$$C�LASS  ����������� VERSION��  �1N�$'  1 ~� T����M-900i�B/700���  �aiS40�/4000 16�0A��
H1 DSP1-S1��	P01.0e�,  	��  ��� � �# ������������
=���r9  w����:��D @m�B  ���� � �t��  ��T��< 7.�7.������ M�  2��'���>U�����\+?��������&Ѡ! ��o�� _���U������= #����I�2�����[�����!B	� � 2 ��� �� �:?���'b�(�/�/�/�/��<?���/A?�S?e?��2�#g���=��<��&��3�V�0��n��W�1�p?�?���0)BT2^2fxk �H��{����@�
(v�F��R�oP�P���^%�  :fd���6}�D�� ���
�	I�)�� ����� e@:"��?�����i\'
���(n����sr'H~/�/��/`q_�_�_�_7а_�>3�_�_oo1oCo�Uogoyoj�?0�?T3^�R"O|BO�TC�lO~Gl�N���y/y/�O  �8� 	��8D�����lU?#�F�O, ���� &8$��zoR$�\,@�����*X� 6_H_Z_#�5�G�Y��-3@h���f���� ŏ׏�����1��o��o aiF/22/3�a8QYe4^4�o�k@Du$������A2���VOZ�&r�� X�$+ ������K>���}#�5�����p��@aq;!�<E�R#J��\!T�����8ߓ�mt&��!y7�@�B ��������	}������4� ���F�k�}�����0��ſ׿�KF�0)j�T5^5����F���8Ɵ؟����������τ����X��c�u� �������R
"�����)(,V3����ʯ�ߥ߷� ��$���H���#�5�G�`Y�k�}������R0"�T6^6FτX�j��s �ϒ��x �n���ϟ�����%�@�p��< �����~������	��� � s�-U^�p߂� K]o��ߐ � ���#5GY������@Z�Ann�	��a����// &/8/J/\/n/�/�/�/ �/�/�/�/�/?"?2<�2?V?h?z?�?�?�?@�?�?�?�?
OC�����EXTE�NDED AXI�S��  T�olmtcGSW�A10����H �a -�����k�C�`���{��q����8��<�AQ�7A� 5�x_
 zD�Hv���O__1_C_��w �[��\��rq!pP��>E��sp�9?
=���5O_�_~�_nQ����`��� ��Bf � 1  
 ����_'o9oKo]o�oo�o�o�o�o�o� ���o���HZ l~������ �� �2�D�V�h�z� ����B?ԏ���
� �.�@�R�d�v�I�o �o��&8 ��$� 6�H�Z�l�~������� Ưد���� �2�D� V���z�������¿Կ ���
��.ϊ����� w�ҟ䟬Ͼ������� ��*�<�N�`�r߄� �ߨߺ��������^� &�8�J�\�n���� ��������H�Z��~� �Ϣ�j�|��������� ������0BT fx������ �,>Pbt ����&���<�N� `�(/:/L/^/p/�/�/ �/�/�/�/�/ ??$? 6?H?Z?l?~?��?�? �?�?�?�?O O2ODO VO����O�/�O �O�O
__._@_R_d_ v_�_�_�_�_�_�_�_ oo*o�?No`oro�o �o�o�o�o�o�o pO�O,�O�O�O�� ������"�4� F�X�j�|�������ď ֏�Do��0�B�T� f�x���������N @�dv�P�b�t� ��������ί��� �(�:�L�^�p����� ���ʿܿ� ��$� 6�H�Z�l�~�ڟ��� ��"�4���� �2�D� V�h�zߌߞ߰����� ����
��.�@�R﮿ v����������� ��*�<��Ϫ�T��� ���Ϻ������� &8J\n��� �����l�4 FXj|���� ��D�v�h�/���� ��x/�/�/�/�/�/�/ �/??,?>?P?b?t? �?�?�?�?�?*�?O O(O:OLO^OpO�O�O �O/8/&/�OJ/\/$_ 6_H_Z_l_~_�_�_�_ �_�_�_�_o o2oDo Vohozo�?�o�o�o�o �o�o
.@Rd �O�O|�O__�� ��*�<�N�`�r��� ������̏ޏ���� &�8��o\�n������� ��ȟڟ����l� �:��������į ֯�����0�B�T� f�x���������ҿ� ��R��,�>�P�b�t� �ϘϪϼ���*�`�N� �r���L�^�p߂ߔ� �߸������� ��$� 6�H�Z�l�~����� ��������� �2�D� V�h�z������Ϥ�� 0�B�
.@Rd v������� *<N`�� ������// &/8/������b/����  �/�/�/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?OOzBOTO fOxO�O�O�O�O�O�O �OR/�/v/?_�/�/t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o&O�o $ 6HZl~��� _"_�F_X_j_2�D� V�h�z�������ԏ ���
��.�@�R�d� v����o����П��� ��*�<�N�`��� �����(���� &�8�J�\�n������� ��ȿڿ����"�4� FϢ�j�|ώϠϲ��� ��������z����� g�¯ԯ�߮������� ����,�>�P�b�t� �����������N� �(�:�L�^�p����� ��������8�J���n� �ߒ�Zl~��� ���� 2D Vhz����� ��
//./@/R/d/ v/�/���/,> P?*?<?N?`?r?�? �?�?�?�?�?�?OO &O8OJO\OnO��O�O �O�O�O�O�O_"_4_ F_�/�/�/�_�/�/�_ �_�_�_oo0oBoTo foxo�o�o�o�o�o�o �ovO>Pbt �������� `_r_��_�_�_���� ����ʏ܏� ��$� 6�H�Z�l�~������� Ɵ؟4��� �2�D� V�h�z��������>� 0�گT�f�x�@�R�d� v���������п��� ��*�<�N�`�rτ� ������������ &�8�J�\�n�ʯ �� ���$������"�4� F�X�j�|������ ��������0�B��� f�x������������� ��,�ߚ�D�� ���ߪ���� (:L^p�� ����� /\�$/ 6/H/Z/l/~/�/�/�/ �/�/4fX?|� �h?z?�?�?�?�?�? �?�?
OO.O@OROdO vO�O�O�O�O/�O�O __*_<_N_`_r_�_ �_�/(??�_:?L?o &o8oJo\ono�o�o�o �o�o�o�o�o"4 FXj�O���� �����0�B�T� �_�_l��_�_
oҏ� ����,�>�P�b�t� ��������Ο���� �(��L�^�p����� ����ʯܯ� �\��� ��*�����ȏ������ ƿؿ���� �2�D� V�h�zόϞϰ����� ��B�
��.�@�R�d� v߈ߚ߬߾��P�>� �b�t�<�N�`�r�� ������������ &�8�J�\�n������� ����������"4 FXj|���ߔ�  �2��0BT fx������ �//,/>/P/��t/ �/�/�/�/�/�/�/? ?(?���R?�� ��?�?�?�? OO$O 6OHOZOlO~O�O�O�O �O�O�O�O_j/2_D_ V_h_z_�_�_�_�_�_ �_B?x?f?/o�?�?do vo�o�o�o�o�o�o�o *<N`r� ���_���� &�8�J�\�n�������  oo��6oHoZo"�4� F�X�j�|�������ğ ֟�����0�B�T� f�x��������ү� ����,�>�P���ޏ Џz������� �(�:�L�^�pςϔ� �ϸ������� ��$� 6ߒ�Z�l�~ߐߢߴ� ���������j����� WﲿĿ�������� ����
��.�@�R�d� v�������������>� *<N`r� ����(�:��^� p��J\n��� �����/"/4/ F/X/j/|/�/�/���/ �/�/�/??0?B?T? f?x?���?. @OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_�/�_�_ �_�_�_�_�_ oo$o 6o�?�?�?o�?�?�o �o�o�o�o 2D Vhz����� ��
�f_.�@�R�d� v���������Џ�� Pobo��o�o�or��� ������̟ޟ��� &�8�J�\�n������� ��ȯ$�����"�4� F�X�j�|�������.�  �ʿD�V�h�0�B�T� f�xϊϜϮ������� ����,�>�P�b�t� ��⯪߼�������� �(�:�L�^ﺿ�޿ �������� ��$� 6�H�Z�l�~������� �������� 2�� Vhz����� ��
x��4�� ��������� //*/</N/`/r/�/ �/�/�/�/�/�/L? &?8?J?\?n?�?�?�? �?�?$VH�?l~ �XOjO|O�O�O�O�O �O�O�O__0_B_T_ f_x_�_�_�_
?�_�_ �_oo,o>oPoboto �o�?OO�o*O<O (:L^p�� ����� ��$� 6�H�Z��_~������� Ə؏���� �2�D� �o�o\��o�o�oԟ ���
��.�@�R�d� v���������Я��� ��t�<�N�`�r��� ������̿޿�L�~� p�ϔ������ϒϤ� �����������"�4� F�X�j�|ߎߠ߲��� ��2�����0�B�T� f�x����
�@�.� ��R�d�,�>�P�b�t� �������������� (:L^p��� ����� $ 6HZl������ �"���/ /2/D/ V/h/z/�/�/�/�/�/ �/�/
??.?@?�d? v?�?�?�?�?�?�?�? OOt��BO�� ��O�O�O�O�O__ &_8_J_\_n_�_�_�_ �_�_�_�_�_Z?"o4o FoXojo|o�o�o�o�o �o2OhOVOzO�OT fx������ ���,�>�P�b�t� ������oΏ���� �(�:�L�^�p����� �o��&8J�$� 6�H�Z�l�~������� Ưد���� �2�D� V�h�ď������¿Կ ���
��.�@Ϝ�Ο ��j����������� ��*�<�N�`�r߄� �ߨߺ��������� &J�\�n���� ����������Zϐ�~� G��ϴ�|��������� ������0BT fx�����.� �,>Pbt �����*��N� `�r�:/L/^/p/�/�/ �/�/�/�/�/ ??$? 6?H?Z?l?~?�?��? �?�?�?�?O O2ODO VOhO����O// 0/�O
__._@_R_d_ v_�_�_�_�_�_�_�_ oo*o<oNo�?ro�o �o�o�o�o�o�o &�O�O�Oo�O�O� ������"�4� F�X�j�|�������ď ֏���Vo�0�B�T� f�x���������ҟ� @R��v��b�t� ��������ί��� �(�:�L�^�p����� �����ܿ� ��$� 6�H�Z�l�~ϐ��� ���4�F�X� �2�D� V�h�zߌߞ߰����� ����
��.�@�R�d� v�ҿ���������� ��*�<�N������� ����������� &8J\n��� �����"~� FXj|���� ���/h�z�$/�� �����/�/�/�/�/�/ �/??,?>?P?b?t? �?�?�?�?�?�?<O O(O:OLO^OpO�O�O �O�O/F/8/�O\/n/ �/H_Z_l_~_�_�_�_ �_�_�_�_o o2oDo Vohozo�o�o�?�o�o �o�o
.@Rd v�O_�O�_,_� ��*�<�N�`�r��� ������̏ޏ���� &�8�J��on������� ��ȟڟ����"�4� ��L������į ֯�����0�B�T� f�x���������ҿ� ���d�,�>�P�b�t� �ϘϪϼ�����<�n� `�
߄�����p߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��"������ �2�D� V�h�z�������0�� ��B�T�.@Rd v������� *<N`r�� ������// &/8/J/\/����t/��  �/�/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0O�TO fOxO�O�O�O�O�O�O �O_d/�/�/2_�/�/ �/�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�oJO$ 6HZl~��� �"_X_F_�j_|_D� V�h�z�������ԏ ���
��.�@�R�d� v������o��П��� ��*�<�N�`�r��� �����(�:��� &�8�J�\�n������� ��ȿڿ����"�4� F�Xϴ�|ώϠϲ��� ��������0ߌ��� ��Z�ԯ��������� ����,�>�P�b�t� ������������ �r�:�L�^�p����� ����������J߀�n� 7�ߤ�l~��� ���� 2D Vhz����� ��
//./@/R/d/ v/�/�/�/�/> Pb*?<?N?`?r?�? �?�?�?�?�?�?OO &O8OJO\OnO�O��O �O�O�O�O�O_"_4_�F_X_�/�$SBR�2 1�%�P� T0 � �C�/�' �_�_�_ �_oo&o8oJo\ono �o�o�o�o�Q�o�_ �o'9K]o �������o� �o#�5�G�Y�k�}��� ����ŏ׏����� 1��U�g�y������� ��ӟ���	��-�?� "�c�F���������ϯ ����)�;�M�_� q�T���x���˿ݿ� ��%�7�I�[�m���ϣφ�~i_� ���� ����*�<�N�`�r߀�ߖߨߺ����ƙQ �Ϡ��#�5�G�Y�k� }������������ ���0�B�T�f�x��� ������������ ,���\n��� �����"4 FX<f���� ���//0/B/T/ f/x/�/n�/�/�/�/ �/??,?>?P?b?t? �?�?�?�?�/�?�?O O(O:OLO^OpO�O�O �O�O�O�O�O�?_$_ 6_H_Z_l_~_�_�_�_ �_�_�_�_o o_Do Vohozo�o�o�o�o�o �o�o
.@R6o v������� ��*�<�N�`�r��� h����̏ޏ���� &�8�J�\�n������� ����ڟ����"�4� F�X�j�|�������į ֯��̟��0�B�T� f�x���������ҿ� �����>�P�b�t� �ϘϪϼ�������� �(�:��^�p߂ߔ� �߸������� ��$� 6�H�Z�l�Pߐ��� ��������� �2�D� V�h�z����������� ����
.@Rd v�������� *<N`r� ������/� &/8/J/\/n/�/�/�/ �/�/�/�/�/?"?4? /X?j?|?�?�?�?�? �?�?�?OO0OBOTO 8?J?�O�O�O�O�O�O �O__,_>_P_b_t_ �_jO|O�_�_�_�_o o(o:oLo^opo�o�o �o�o�_�o�o $ 6HZl~��� ����o� �2�D� V�h�z�������ԏ ���
�� �@�R�d� v���������П��� ��*�<�N�2�r��� ������̯ޯ��� &�8�J�\�n���d��� ��ȿڿ����"�4� F�X�j�|ώϠϲϖ� ��������0�B�T� f�xߊߜ߮������� ����,�>�P�b�t� ������������ ����:�L�^�p����� ���������� $ 6�,�l~��� ���� 2D VhLv���� ��
//./@/R/d/ v/�/�/~�/�/�/�/ ??*?<?N?`?r?�? �?�?�?�?�/�?OO &O8OJO\OnO�O�O�O �O�O�O�O�O�?"_4_ F_X_j_|_�_�_�_�_ �_�_�_oo0o_To foxo�o�o�o�o�o�o �o,>PbFo �������� �(�:�L�^�p����� x��ʏ܏� ��$� 6�H�Z�l�~������� �������� �2�D� V�h�z�������¯ԯ �ʟܟ�.�@�R�d� v���������п��� ����&�N�`�rτ� �ϨϺ��������� &�8�J�.�n߀ߒߤ� �����������"�4� F�X�j�|�`ߠ���� ��������0�B�T� f�x������������� ��,>Pbt �������� (:L^p�� ����� //� 6/H/Z/l/~/�/�/�/ �/�/�/�/? ?2?D? (/h?z?�?�?�?�?�? �?�?
OO.O@OROdO H?Z?�O�O�O�O�O�O __*_<_N_`_r_�_ �_zO�O�_�_�_oo &o8oJo\ono�o�o�o �o�o�_�o�o"4 FXj|���� ����o�0�B�T� f�x���������ҏ� ����,��P�b�t� ��������Ο���� �(�:�L�^�B����� ����ʯܯ� ��$� 6�H�Z�l�~���t��� ƿؿ���� �2�D� V�h�zόϞϰ��Ϧ� ����
��.�@�R�d� v߈ߚ߬߾������� ���*�<�N�`�r�� ������������ ��
�J�\�n������� ����������"4 F*�<�|���� ���0BT fx\����� �//,/>/P/b/t/ �/�/�/��/�/�/? ?(?:?L?^?p?�?�? �?�?�?�?�/ OO$O 6OHOZOlO~O�O�O�O �O�O�O�O_�?2_D_ V_h_z_�_�_�_�_�_ �_�_
oo.o@o$_do vo�o�o�o�o�o�o�o *<N`rVo �������� &�8�J�\�n������� �ȏڏ����"�4� F�X�j�|�������ğ ��������0�B�T� f�x���������ү� ��ڟ�,�>�P�b�t� ��������ο��� �(��6�^�pςϔ� �ϸ������� ��$� 6�H�Z�>�~ߐߢߴ� ��������� �2�D� V�h�z��p߰����� ����
��.�@�R�d� v��������������� *<N`r� �������� &8J\n��� �����/"/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? 8/x?�?�?�?�?�?�? �?OO,O>OPObOtO X?j?�O�O�O�O�O_ _(_:_L_^_p_�_�_ �_�O�O�_�_ oo$o 6oHoZolo~o�o�o�o �o�o�_�o 2D Vhz����� ��
��o.�@�R�d� v���������Џ�� ��*�<�N�