��   A��A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ������DMR_S�HFERR_T �  $O�FFSET  � 	4/GR�P: $�MA��R_DON�E  $OT�_MINUSJ � 	sPLzdC�OUNJ$REF,j�PO{���I$BCKLSH�_SIG�EA�CHMSTj�SsPC�
�MOVn �~ADAPT_I�NERJ FR�ICCOL_Pz,MGRAV��� HISID�SPk�HIFT�_7 O �N\m�MCH� S��ARM_PARA�O dcANG�o y2�CLD�E7�CALIB�Dn$GEA�R�2(��� RING��<�$]_d�REL�3� 1  	��P CLo: �� �AX{  �$PS_�TI����TIME ��J� _CMD,��"FB�VS �&�CL_OV�� F�RMZ�$DED�X�$NA� %��CURL�W����TCK5�wFMSV�M_LIF	��`;8G:w$�A9_0M:_��=�93x6W� |�"�PCCOM���FB� M�0�M7AL_�ECIr�PL!�"DTYk�R_�"�5L#�1EN�DD��o1� �5M�P PL|� W �  $�STAL#TRQ_�M��0KN}FSD� �HY�J� |GI�JeI�JI�E#3AnC�uB�A�4�$�A{SS> ���	Q������@VER�SI� W  1N�$S� 1'X ���� 	 ���n_Y_�_}V*v� ix x,���� F���\m���XZ6�?8�6��G�_S���8��G����P��P��l��#m�u_� *k�S�oQTo�]�J���I\ �������oh��$b�Ao�o�_gl�o �o�ot� 7uޗg@Mv @
BZpYq#�o�su���Ef ��ZVPm
P�  k��dw������=L���.�?�/���@�O�t��� ������Ώ�����(�:�� 	Ue�s�8]���T  2�ğ ֟�����0�B�T�f��R��������Ư د���� �2�D�V� h�z�������¿Կ� ��
��.�@�R�d�v� �ϚϬϾ�������� �*�<�N�`�r߄ߖ� �ߺ���������&� 8�J�\�n������<���������&��8�J�\�n������|( u��q������2 /hS�w�� ���
U_.�R=�K�5`I �E�o��/s���,///T/z/��/�/�/�/�/�#�<h/f C@�/*? e/N?9?r?�y���?�? �?�?�?�?OO/OAO SOeOwO�O���O�O�O �O�O_R��Ov�(_^_ ���_�_�_�_�_�_�_ oo'or�Ko]ooo�o �o�o�o�o�o�o�o #5GYk}�� �������1� C�U�g�y��������� ӏ���	��-�?�Q� c�u���������ϟ� ���)�;�M�_��� Ho������˯ݯ�� �%�7�I�[������� d?����ٿĿ���!� 3��W�B�{�fϟϊ����s��$FMS_�GRP 1mU� ����P\R�J����J���N���K1UIM�����GC@uM���M���H��JJ�nKG�r���A�V߯���.�A�@h��6�&;�w�1c{BX�/�π�߭�T�fߠ���R����/��S�>��w��R� 6�S]bn�r�� � �����z�B�A�L���6E�;*�1��BY*tn��G�A���6�2�:L�\�1��2BY;3b�>��T@B&�����Y���)>����Js��2  }  ��%CC_AU�T01��s��x� tS����������� }�Z�+~���a��� p�� �D� 'K6o��� �
�V�/�5/ G/�k/���//�/ �/�/�/N/`/1?�/�/ g?R?�?v?�?�??�? 8?J?O�?OQO<OuO �O�?�O�?O�O\O_ �O_;_�O�Oq_�O&_ �_�_�_�_�_oT_%o x_�_[o�_Xo�o|o�o �oo�o>oPo!�oE 0U{�o�o�f ����/�A��e� �������я���� �Z�+�~���a�܏�� p������ ��D��� '��K�6�o���ԟ�� ��
�ۯV�د���5� G���k���Я���ſ ��տ��N�`�1τ�� g�Rϋ�vϯ������ 8�J�ߖ��Q�<�u�����ϫ���g�4� ����[���W���2��<V�A��P{]�`��������I�RG� ���#���)��,�Q�w� �_��y��� � ��R�"����󙚭�T��N<����@Q��	���  ���TOD_GU��f>��������ѿzy�g�/�����	J|���d�F ��not �a progra�m�.����'�8yZ��)�ad�)"��t�|
���*�D����+�b!/$/���I/����/6|	2#~��/L/��,�x�/�/���	?t/�/�/i?�*�JM`q??�(�J�?�?�+�B��?4?F?X?)O|	 �����81O�?�*si�aOdO:�@�O�OD�O�O�O� _X�9_$_I_o_��O �_s_�_O_�_�_�_ .o�_�_do�_o�oo �o�o�o�oGoko}o N`K�o�� �1C��8�#�5� n������Y�ڏU� ���"�4���X����� ������ğ�����M� �q���T�ϟx�c�u� �����7������ >�)�b�t�ǯ����� ο�˿��(�:ύ� ^ϱ�ÿ��ϸϣϵ� ��A�S�$�w���Z��� ~�iߢߴ����+�=� � ��D�/�h�z��������[�����$P�LCL_GRP �1������� p�>���?�  �x?XS?r����� E���i�T���x����� ��������/6K������r�5?}"�(�!��# ����� 2 VAze��� 