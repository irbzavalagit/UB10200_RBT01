��   ��A��*SYST�EM*��V9.3�0126 2/�12/2021 �A ��������TW_CAPC�FG_T   �\$MAXW�EAR_FIX w BMOVNALARMSE]�$RESERV�EDkIOTYP�xIDM$SA�V_DATEN �/PRM6 ��$MINWR�4CALC^p
S?TD_VALJK �_TOL_NEG�
POSN�[[ ��
}�4/M�EAS9 �$_Iw_CT��TIPqSPOT|_=p
3 FK��[COMPp Sp��[FRATK��PC� ��_IO_OBC�S�<%�_."NZ�AV8 l��ED�ABL�E�%�1~2�N�UM_TE� �T�IMESTAMP!�'�!�� T2~9 0$� �U��$~|�$���ZGUN9�@ '�6  	 �?3%N5�]6�=$N5=0HI� IM��"�4|�4FF_4�DIF�p�#PL�S_ZRO�"$O�PN� �"Q `B0ƗME�0�0FEN	Do B0�I E`�,F=$I@MX� SG� `D!\HvB lG!!\H�BlC<"C ]C�E�HvH�G�DALI�B�$EXTRA_INT�#�F�3�C/REAL�!X�3���1�1w<WK W�Y >SYX$4��6� � �4�0RQ�3S_�1V� ��3�Q�3� �3ENBL�N + QCHMS��$DRAM_�FLOORQSRO|�Y�P_MASK�O�__*Y4�$$�CLASS  O���Oa��`���`D`VERSIO�NLh  1N�$TW+0y100mh`A ��4�`Ub��?��d��X�d�j�lBH����c0�i�e��e@�sz��h%7 hJr ��MF���Aߤ  �` ��?�`>o���p:�`�qA���Bi��B&V.OaRru��``p�`fq�>L� >!��ruA>���`fM��B)�l�~�� �d���
����jq�aSQ�nqR�2��w���������R��,���bx`��~eV1�  �jJp ;�s��0�`Q����
�2:�� ��
�\��*"
�3��c�4���a�
�5ß՜6� �Q�
�7� SE
�8)�bq
�9K�L�2�o�o�o�o�o�o �o.�:I�d�v� ��������п���� �*�<�N�`�rτϖ� �Ϻ����υ��Ӝ�����.�����/�~��c߲�-�2������5��/��/�(�`�J���l���~d3������ïկ��� ��5�A�P�k�}��� ������������ 1CUgy��� ������ϱ�� ߀��j/�3�ߝ��ԛ3��X� /�Q�sﲘzS �P~,hp�s��c���