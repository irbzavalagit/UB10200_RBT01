��   4��A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ����SG_LOG�ARR_T� �$CLK  �$MCHPOS�= $CMDET�RQ= $HPD�^DTMAXfI�N^FCSTAT�zMeERROR�_CNT3=XT�RA_SHORT�1^�2���	4�^�4&CFG�0 � $G�UN_NUM_M�S<CURFNO4ROO�m * �_OPT�&DB�G/�INTVA�RGFRELOF�ILWRTTMM�o* STRTWTsLMC* TYPRPS_�L��L��\������&INF0, &'�=��=SG(�$A�CTVRQSTC�Oe . IDoT�RKIDK- fA�T� MP="$�TMH+OTLl C�C"�Nkk&TA�SK$$� RT�RE ?$OSTI�ME=ROUT_�N��$�#COwMME�%'�hAB� ^RESERVED�* t!;_T�PRS)0m )_DU?#�0LONG�21�21P�21�:857;67;77;8�A��1� �7��8��8r1�8�1��8�1�8�1�h0� �7 � �gIG!�<C5#ALINC���%��)�E%hP)�EhSAV_EPATHP %�ENA�!� -??>�?���0� �(�%�� (ENB= 'TRI6�.��'USE_??��MDEST_DI�R%RhNM_BAcSE�V�nINz�N�� YS_FL=GUFFORM���EVT� x �
�!TUG$T�]D�AN�Q�PA�PCLOC<*-%�SPEEeTHI_CKNESGE�F\=bcFLO���� �� 2$�WELD�`Ze�_�TO\CONT_�SdCLSTHRS�@Qb�`��b��b���c�fDST1qC�P�c�PST2y��OBRk+xAV�*-r�PTj #PDbRsYq6wcsINky�Dy,p_TH3PROTsckrk�OM?wb�8dwb�3E�@� 2	`�PXE �."`UjF�CTL_SWIT�C�cP183UN�CLMd6�<�^@E�&E--%PSCHn�&WLDn�SDX�TSK�FLAx�S�T�VCTRLK�HI0Q�OK_M�MHu�`LDDIS��s�'%TCPX_GAF_z�H��Y��UZ��W��P��R���4�$9 A[` O���[���o��moP�VE�`ONX��  1�N�	#AR2 2� [�f� A$[�[�������3��h����ʘR֟ $���=���� � y�o � � cn���'� !>����A#]����b�������������  %�&�ݪ �J�\�n� _�ݢ̯���ſ���\����MEM���t� ��Я���ο�Ϯ�<� �����τ�Gύ�>߉��O�t߆ߒ�� 1  $�~�i���������	�˕��2�߷�,�>�����3	���t������IN2�[���A�'�e� w�Q�5�Z���{�����]���3������a�� )�;�B_�q�u��"��F��e�4���@�;B&Ppt���T 2ٙ�|�%
SPOT?[] log�O***��2�TP�`OT�,v�c� %}�b_MOTN�(��, PN!��,;#B"
΀*�R/^/p/�/�!O�K�+<;#B#Ac�celtime �tun�/�/x?c:TYU�*b�]pF$�
w�C!P113�(dyn fri?ction)Q?l?��1O�?�$�0�<�5�P47(inertia�?�?���?O�%$H@�?�683(c�losP0hres�hSOkO�O�O!J83�A�O�G�C fct�l2�O�O�_!\B1]�#6�9�JX_k_��_�_![9�Hb��5�6�1(sprin�g consta�nt�_�_oo$X1�0O�V2(p�@su?re gai�?�1�oo?�o%W2�L�%~��2 parm�QP`����o %FC2PARM3�E@Auto Ze�ro calibrateu�o$?AUTOMAW��x���ZDefle��2����-DFL_CTCAL )D����ZManual� �f(gunke�y)�+n���3MA�NPR��1MP�"�UȄweld��/��=�ANWL�DvI*�W"?%P �eS�O�T�n�ӆ�����PC��@$�Tipwear �mea�ament�ܟ���%IPWE�AR�T���%P�oke schedule[�g�y��OKRE�J*����5:A3ȢtesZ��s��� TS/**�/+�;a?5MoN�ev�̀R�f���MOkEV��@>h�anel sL�c�hП��oO�O"SR#CH�����>HI�detL�Կj�|ώ'PANELDE%�߽�ȖChe�ck����ʇ��HH7����(�P Π T�bt߆ϬQ�����Ac	Reserved1�c��߇][�����G�(��m������G�3������0�]���=�d4Y���`u�������d5�c���]�=d6�Ycu��d7��]���XtraP���p���!XTRA��"_�  ��$SG��IN2 �2'�S!o� /t/�/ �S!�%�)�� �/�/ �/�/??'?9?K?]? o?�?�?�?�?�?�?�?�+MU#%/6O�/�' dOvO�O�/�/�O�O�O �O__*_<_N_`_r_ �_�_�_�_�_�_�_O O&o8oKO]Ono�o�O Io�O�o�o�o�o" 4FXj|��� ����ooo0�Co�lF&3P/b/�����o �o������!�3�E� W�i�{�������ß՟ ���� ��$�S� Zo����Z���ҏ��� ��+�=�O�a�s��� ������Ϳ߿��� (�:�K�^�l�Xϓϥ� ��ʯ�������#�5� G�Y�k�}ߏߡ߳��� ������� �2��U����\�Fn� D�j��& ?�����X�����,���� e��������'� � ������)�$#�r�p��J��V�'� �R�%���p�0��V�&�~�������*�@穙���� W�� 2� '%	S012SSW0��)E��Z��Æ|�=������C@0z/v������� /ASew�� �����//+/  �2�6/s/�zϩ/�/ z/�/�??'?9?K? ]?o?�?�?�?�?�?�? �?�?O#O5OH/Z/kO ~/�M