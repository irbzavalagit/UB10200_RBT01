��   	s�A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ����SG_BAC�KUP_T  � ( $COM�MENT �$STROKE � $USE_�MANUALL �4�$$CLAS�S  ����k����` VE�RSIONh�  1N��$SG*1 1 ��u 	G�un Close���	10mm_ Open�� �U2���3����	4�
B�5�H�6p7��8�9��
10�	Bm��
1�
Bܡ��
B
1C̡C�1C��IC(
1aC���yC4��C>�2�C@�!�
3CR�&�
C\�&��f�&
+X
2"+z$�&:+��&R+��&j+�p
2�+���2 ������! 3EWi{��� ����////A/ S/e/w/�/�/�/�/�/ �/�/??+?=?O?a?s?�73�?�0���3�o �o�o�o�o�o�o' 4FXo|��� ������0�G� T�f�x���������׏ �����,�U�