��   �6�A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ����SW_ADV�FUNC_T �  P $FA�STFLTREC�  $AUT�O_REWELD�ENUMN TRI[ESE $^YN �GeMOTION�_LOCKE4�&CELL1 �L8 HOME_P�OS_PReSHގPOLLEPB�_NOQ�STR�OKE�SOPR�UNE�IO1�t 7$DO_�JTe�IMA�NUA�PR�CALT 8CLRXFR XOPENCx�REP|�ATPNCE ������/? >�N�OTAB�$W�DENB4$/COM>W!��7*t$�PRTI��#��RQ   8�(�&MNT�,�#>�(OUTTO�,��(IWV+ 4I_�LV� >576RT�HMF�\6U7PC�MP|6U7MTW1S]�6�:LD�;�0��9� �:�1k'IMI�NFz(�3�=� ��1SP=.B'DaX� (KC�#
·�ONFIG1�< &YWD_C�TLS ��_�6!EQ�GLCH_�FFe 0_TYP�E�BTD_AFT�ER_CD�@DU_MP_CH�$�0_HID��A�F�A�CYCLc�ADE9FZ 	VWDU��A�VENDO�$�PS�@_DSB_-D��$<UE�A�@�TDFFEXCH�ri �BPREV<ERCOUNXP�N C_O�GWAR~�$CUSTOS�o@T�A�@�WOND�LY�XF�UFRCΝ1NWDH LR�\ CVRS�@I��@SP�AeEXT�_WSD_SCH~UDX_CFG� �PdA$OK2SK�P_SPO�S�QC�NF�FQWKVI�EWd�BSHRTFTnIT�SJ�0IT�SNlPLOaS`TwRNSfZDT7�Te�EQ� { ^T_GUN�)�d�(STtA�j�(|#BU�lp�(Q~2t�)P|Vs�(�4py�(#HV��y�(M�{�q��(@0�)�q�%GO_?BINMPV�&�w �y���y�2��y�P��{EQ7k��(�`aC�P�(���yD1:ං��zւmz_BY9P��*OB�y5!8^9�ODER]W��`PRS��w��(��;����:��/EN�W=ْ76WSOK��'���&��F���MW_FLW
�6����C�`Sy�X�����I����VC\��2�����X�Ƣ��BUOP����۪C�3 ���G�	�*����J���TC�GN�P�p�e�NESQ�����H^ 
������AIR�3һ��HD�h���x���yE78�76NS�Põ?(�?�?�=G6�A� q�x���dSETU�?p IY�`.TTUDQE�VQUDBACKU�Q�VRDROPO�A�%WQPI ���2x�0ӟBCTRL����#G_SEQUE#NT��a��Rd� �RE^��AfPULdS��PTa{`NT4�1OT�PrB4���a��o�� T_�UVp�a��@��p��p _ID�X�$SOF=OU�a ���Ѯ@TI Sp��q|��ӻ�x�P��6�DELA�S�v�G�QU�WOS. �WCU�cOo�$q�MUL��u��Z`��![���EQ�P:��Vt@MB4w�c,r���AF��P�@s {AT.�EPB4� G�S�A@!��EV)�C���E I*�c�D��pC�  #�|�"|�x!�Vp ��g҃�����l�T  �����R��jQ��` �GGN���OO�@G �abS����g����G�J�B{��Ü�FT��}xGN|PEuD��A�CCLS�cEM��L�0�uE�N�@ ��`M� O�R ��O�I�Q��A%c~t�OC_NAMn��	$/Po�4PA�U�����uA ,K �CO��!L"]F" DP�4a�_TS� D~+STYLE_S���CE�XTRA_SHORT1&�]Q�_MS�A������ßA�c�� �$MAJORb�@Gc @�EO;��|ּ�$A�%SS T�l֭RE+Po@|�P�D0IME�S"M_3FA�AR�ST�AF̂"PST`�PMEDLA��D��o�#0��$Iv�DLVL�"#ARL `�cHT�o���K+@>T%$ARITYz�+@9 p��%:���`CHE��I5k�o�Pr`3Fi4��D�!���3`79�OH�4�7Tw�ܘ�4���#�;>k�USER12GC
�:2K2�9��HCDp:K)HcD�7EFEN3����C�����9}9FW��#�Lk�MDSONT��F�ITW��Kk��ALH��%Tk�OP�KET�7Hl��HeTM�CAP5\��S�7Qu��8�Sk�E���X�Tk�INRQT;��Z�8�INIn9ck�WD����4� g���5KCH�?jB6�O8ed� +;�f�`�!�l�h�I��f�h�9�f��AL1Mr�t�gIN{&s ��!FCu<z)Fau�iP(Gv햅AIx�s�z8gx�s�CFL�h�s`�{�y�s�6�AR
x<��AHDBg�s�D;��M�i[��hI�i{�|gOTO�h����AUT
V���CROV��Մ��i2�U�c�k0�W�<wAu�Q@Jx6�,��XS��T�p89�u�|gNRD�W�����pCO�ȵ�d��|��7$LEA�� ��+d��:f�K��"�<��DEV_N��+d8 ��"&NDX��t @��(0@�(ZS��C
N�T�s�j�WC���dܘ��4��_B�N� 	 X ��4CЬ��D?UR10TH����DOSf!O������CF�Q
 H`+�H`�0�AL��SEV�ĢD��MSG�c�Հ|�[TM��$��A��� ��%���ڇ� ��VE�RSIe���  1N�$��ADVFUNC�  ������ݶ����C?ELL ��׶2ܹ�~���رD��:�47�Y�k�3g̭1g��g�2gĵ*i�g��ı=Ī���ϩ�ݵj�ܵ�ϸ��ܱ��ܱ�� S�im infor+m:�˽g�
��]��ݸ�ONFIG �̿�ܹƏ�� ˰�߱��ߙ�P�5 ����ܱ豚��OOM  ��װ�������k̡�lߌEQv%�1����� k�������,�>������B�T�~�������������������B ����9K]o��i���*�k�
�� �� 2DVhz �������
/�/./@/R/��/�� ���/�/�/�/�/? ?/?A?S?_?q?�? �?w?�?�?�?OO+O =O����Fd/�O �O�O�O�O__0_B_ T_f_x_�_�_�_�_�_ �_�_oo�ONo�/JO to�o�o�o�o�o�o�o �?�?4^p� L����� ��O tO&�Xo�O0o6o���� ��Ə؏���� �2� D�V�h�z������� ԟ�`��lo�@�R� d�v���������Я� �� �*�<�N��Z� ��������̿.�@�� d�v����\�nπϒ� �϶����������"� 4�F�X�j�|ߎߠ�� �&�����0�B� T�f�x����p��� ���������&�P�b� t����������0Ϧ� T�
(:L^p� ������  $6HZl�������$SPOTEQ�SETUP 1������ ��� %$*�
.�-//@Q/</u/`+��+ȶE,A�*����} �*�!�/?!?3?8������$�8�9��A�  @@D?  Ж2�?�?�?A?h�?���C�/T�?A�d>D
B��JC M��	a0�� �Oa/�O�O�O�O�O_ �/�/�/�/�/�?�/�? �_�_�_��`;�bv: 0�_�?*o<oNolo.O OO�o:LA�MO�oqO �O,�OP;M�q �%_�oI_�om_o�_ �A�S�e��_�_oQo coŏ׏y���o�o�o ��o�o�oƟ� �՟� ��D��� ����+��ۯ� �����������_�q� ���'�9�g���o��� ������`�+���oϨ� �ϥ���Y�k�}����� #�ů��u߇ߙ��1� C���������;��� ӿ�S�	��-Ϛ��TAT 1� ��<����	���!�� h�?�����u���������������NUME�Q  �����S0ALARM9_0�H�S0CLOSEZ~lCHMIN1{��TSKINFO� 2��  ��`1��`0M���	�);M_ q��������//���WELD�IO 1�� 
���Y�;�(�O2��� q$�n�g!��q'Dŋ"O3��� A��(�(��$��$� �/�,+Ӱ!5��/*?<?N?�!��,ĵ$�-E�VE���44��4��4��;�?�?�?O�OJ�!Ot!�1�:�4�-M
0oF9O
�:[2
�O@ȞO �O?˩�[*�s/�+(� �/�?V?t_�_�_?? �_�_�_oV_ o�OLo ^opo�o�o�o�o�o8O �o�nmO�o�ON`�O �g�O_!_3_E_/o o�1�C��_�_y��� �����ˏ1��	�� -�?�Q�c�u��o���� ��=���s0�� �����ۏŏ˯ ݯ�]�o�%�7�I�[� ��w�ݟ����ǿٿ� ���!Ϗ�E�/�şS� 韦ϸ���Ͽ�U�g� y�������q�w߉ߛ� 	���������Y�#� ��O�a�s����� ��;�����q����R� d��ψ�k���%�7� I�3��#5G���� }����5�� 1CUgy�� ����A��/w� 4//����������� ��/�/�/as)?;? M?_?�/{?��?�?�? �?�?OO%O�IO3O �WO��O�O#/�O�O Y/k/}/�/�/�?u?{_ �_�_??�_�_�_o ]_'o�OSoeowo�o�o �o�o�o?O�o�ouO �OVh�O�o__ )_;_M_7o!o'�9�K� �_�_��������	�ӏ 9���#�5�G�Y�k� }��o����!��E� �{8������ ��͏ӯ���e�w� -�?�Q�c����埫� ��Ͽ����)ϗ� M�7�͟[�����'������]��$WLD�CTBNCHMK 2	���!�����4%  *5� <�F��� 2�h�z�Yߞ߰ߏ��� ����
����@�R�1� v��g�������� �����<�N�-�r��� c������������� &J\;��q �����" FX7|�m�� ����/0//T/ f/E/�/i/�/�/�/�/ �/�/?,??P?b?A? �?�?w?�?�����? �?�?�?'OOO]O<O NO�OrO�O�O�O�O�O �O#_5__Y_8_J_�_ n_�_�_�_�_�_�_�_ 1oo"ogoFo�o�o|o �o�o�o�o	�o- cBT�x�� �����;��_� q�P�������ˏݏ�� ����7��(�m�L� ^�������ٟ��ʟ� �3�E�$�i�{�Z��� ����կ��Ư���� A� �2�w�V�h����� ���¿����=�O� .�sυ�dϩψϚ��� ��������K�*�<� ��`�r߷ߖ������� �#��G�Y�8�}�\� n����������� ���U�4�F���j��� ����������- Q0B�fx�� ����)_ >��t���� /�%///[/:/L/ �/p/�/�/�/�/�/�/ �/3??W?i?H?�?�? ~?�?�?�?�?�?�?/O O OeODOVO�OzO�O �O�O�O_�O+_=__ a_s_R_�_�_�_�_�_ �_o�_�_9oo*ooo No`o�o�o�o�o�o�o �o5G&k}\ �������� �C�"�4�y�X�j��� ��ӏ�ď	����?� Q�0�u�T�f������� ���ҟ����M�,� >���b�������ݯ� ί�%��I�(�:�� ^�p��������ʿܿ !� ��W�6�{ύ�l� ���Ϣ���������� �S�2�D߉�h�z߿� �߰�������+�
�O� a�@���v����� ������'���]�<� N���r�������������#5[
�D�aJ�
SGq`~�
�����
��_�+
�z=_
`q�N�
UV���
���
���//
��qo/c/
X�R/�/
�eY�/�/
�ob�/�/
qZ�/3?
��"?g?
�h6V?�?
ǉ��?�?
�8�OT���?7O��+F&OkO
�/q�ZO�O
OxO�O�O
o.�O_���O;_
���*_o_
<�^_�_
����_�_
�E1��_o
^>o�/  .oso
��PPbo�o
�?��o�o
_XE<��oC
�ʏ2w>��f�
��<Ϛ�
��8-o�� ��G�bl6�{�
�?ao��E1+���
ǖ(7ҏ��{���K�
��,`<���Ƥ	�Gn���
6�*���
oP/�ǆ��
�O�
�H8�����
r����
�GN���N[UqMگ�
!!��S�&�$B���
a#]�v���b��YO���޿#�
�qI��V� ��Fό��
&m��υl�Į���R�o&�8��\ߣ
TIߎߠ�� �ߣߵ�������0�� !�f�E�W��{����  �4�����ִ�-�����a�s��R������������� ����9*oN``���� _|���$WLDCTC�FG 
��}��32� 