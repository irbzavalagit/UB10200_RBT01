��   L�A��*SYST�EM*��V9.3�0126 2/�12/2021 A 
  ����CELLSE�T_T  � w$GI_ST�YSEL_P �7T  
7ISO:iRibDiTRA�R|��I_INI; �����bU9A�RTaRSRPNSS1Q23U4567y8Q
TROBQ?ACKSNO� �)�7�E� S�a�o�z�2 3 4 5* 6 7 8aw.n&GINm'D�&� �)%��)4%��)P%���)l%SN�{(O�U��!7� OPT�NA�73�73.:BP<;}a6.:C<;CK;�CaI_DECS�NA�3R�3�TR�Y1��4��4�PTHCN�8D�D>�INCYC@HG��KD�TASKOK�{D�{D�7:�E �U:�Ch6�E�J�6�C�6U�J�6O�;0U��:IATL0RHaRbH<aRBGSOLA�6�VbG�S�MAx��Vp��Tb@SEGq��T��T�@REQ �d�drG�:Mf�G�JO_HFAUL��Xd�dvgALE@� �g�c�g�cvgE� x�H�dvgNDBR�H<�dgRGAB�Xt�b�4�CLM�LIy@   $TYPES�INDEXS�$�$CLASS  ����lq�����apVERSI�ONix ? 1N�$'61j�r���p��q̛t+ UP0 �x�Style �Select 	�  ��r�uReq. /Echo���yAck�s��sInitiat(�p�r�s�t@�O��a�p���	��  U�����������q�������q���sOption? bit A��p��B����C�Dewcis�cod;���zTryout �mL��"Pa�th segJ�n�tin.�II�y�c:��#\�ask� OK��!�Man�ual opt.%r�pAԖBޟԖ�C�� decsn� ِ�Robot� interlo��"�>� isol3��C��i/�"�z�ment��z�ِ���"�^�statu�s�"	MH ?Fault:��'��Aler�#���r�0�p@r 1�z� L��W�i�{���$; LE_COM�NT ?�y� � ��䆳�Ŀֿ �����0�B�T�g� xϊϜϮ��������� ��,�>�P�b�t߆� �ߪ߼��������� (�:�L�����Y����ﾃSY�������p��)���H.S5��G� ��]�o�  �@������0�  ������w� %# I[m���� ���!3EW�i���  x ���H����/� $/J/4/Z/�/j/|/�/ �/�/�/�/�/?4??�0?V?|?f?�?�?t�qȽ>UM�?p�?1�?���?TMOO $O R��ZAIN�NT4OOL\O �$�NMPF�NTR�_�NIF�O�O  �AC�OPTG�OD�_"_  LApOT�NUa_[O $UN��O_P�^CRHOzX��_�?o#o5oGo Yoko}o�o�o�o�o�oP�o�o���-, *dv����� ����*�<�N�`��r���������̏y����	��-���=� c�u������������� А�����/�A�S� e���韛�����ѯ������>�=�O�  (����������� ��ҿ�����,�>πP�b�tφϘϪϼ��Tool Change�������"��4�F�X�j�  yT� Maint�enance P�ospQTip ?Dress ��oR�Reset S?tepper�Ѩ��CC Auto/�ManualoR�Purge Gu'n 1^���2^�\���(�:�L�] D ]�o������� ��&�%�7�I�[�m��W��2@YLE_CO�UNT����������ENAB�  ~����� ����%7 I[m���� ���!3EW i{������ �////A/S/e/w/ �/�/�/�/�/�/�/? ?+?=?O?a?s?�?�?��?�?��E_MEN�U������NA�ME ?%��(%�*D  %O.E  OSO>OwObOtO�O �O�O�O�O�O__=_ (_:_L_^_p_�_�_�_ �_�_�_�_ oo$o]o Ho�olo�o�o�o�o�o �o�o#G2DV hz������ �
��.�@�R���v� ��������Џ��$� ~��S�>�w�b����� ������������=� (�:�L�^��������� ߯ʯ�� ��$�]� H���l���������ƿ ���#��G�2�P�V� h�zό��ϰ������ ��
��.�g�Rߋ�v� �ߚ߸߾�������-� �Q�<�u�`�r��� ��������� �&� 8�J�\����������� ��������7"[F j������ �!E0BTf �������� //,/e/P/�/t/�/ �/�/�/�/?�/+?? O?:?X?^?p?�?�?�? �?�?�?O OO$O6O oOZO�O~O�O�O�O�F甕��O_ �1y�O3_ h=1"_�[_ YOJ_�_ �c�r_�_ �y��_�_ P�P�_��_ LIC�_#o ��oKo  AyG:oso ��bo��o �>�o�o ��W߲o�o јy��o �O��;  �*c ���R� ?�9Qz� n��O��  �y�� �@��+� ��y��S� ASB��{� ?�?j��� �I_Ē�ˏ oy���� ^_p���  �B�  �_ o2�k� oYyZ��� �������� ����� �F�A�
�  ��<1�2�  ���oZ��  �H�J��� � �r��� �y���ӯ ?J¯���  �O�#� � @�K� ��q_r���/[b��� �L���ÿ O����}�KY�ϭ`�|��:�  ��*Ϟc� ;�MRϋ� #��!���%p�)�ϟ  �=���� �� ���+� �y��S� ��Bߞ{� l�jߣ� �_���� �y#���� ����� a!)�B�  �p_i�j�  2�9�Z�� ITyϺ�  M����e�Z�A�����I��3� ����"�[� ��9�J��� VLI_�����S5���� !|I���  NNL���# S��K �IUB:s e9�b� S�џ��  ���� �D@�� @9; �6��b  ��DR��Op����[,d�/ ��q�*/�N/`9/K/]/o/�2��/ �//�/�/�/�/?r�0?i?�&	��?-��?�)?�?�7GRٿ
O � �Sh�?3O �k("O[O�?OjO�ON�DE�O�OO�O�O� ___*_<_Q^CR��O�_5��_Y_�_�Wz��_o�_5o o2oDl�TCHANGE_S221hoJo�o�o �o�l��o&#6yB{>���~�z
MAINT�`�30��xTIPDRESS�q�o���E�rW0B��sC7AP_}f33H��sPURGE1�q�4p��xSTYLE235����ԏ ���1��U�@�R�d��v�����ӟ ��� ������4�J��	:�s������������ʯܯP� �:��� ^�I�[�m������ܿ 7�