��   �A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ����FSAC_L�ST_T   �8 $CLNT�_NAME �!$IP_ADD�RESSB $A�CCN _LVL  $APPP � 4�$8 A~O  ���z�����o VER�SIONw�  1N�$'DEF\ w { ��� ���ENOABLEw ������LIST 2� �  @�!���17�2.19.89.251 Y
��  ��
[ K��H�l~�� ��/��M/ /q/ D/�/h/z/�/�/�/�/ ?�/�/
?[?.?@?�? d?�?�?�?�?�?O�? 3OOWO*O<O�O`O�O �O�O�O�O�O�O__ S_&_8_J_�_n_�_�_�_�_��