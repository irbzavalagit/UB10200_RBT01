��   #��A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG4��DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S?ETHOST���NSS* 8��D�FACE_�NUM? $DBG_LEVEL��OM_NAM� �!�* D �$PRIMAR�_IG !$AL�TERN1�<W?AIT_TIA �� FT� =@� LOG_8	��CMO>$DN�LD_FI:�S�UBDIRCAPΌ �8 . �4� H�ADD�RTYP�H N�GTH��4��z +LS�&�$ROBOT2P�EER2� MAS�K4MRU~OM�GDEV��PI�NFO�  �$$$X4��RCMT �A$| ��QSI�Z�X�� TAT�USWMAILS�ERV $PL�AN� <$LI}N<$CLU����<$TO�P$�CC�&FR�&�J�EC�!�%ENB{ � ALAR�!�B�TP�/3�V�8 S��$VAR79M ON,6��,6oAPPL,6PA� 8-5B +7POR��#�_12ALERT��&�2URL }}�3ATTAC���0ERR_THRO�3US�9�!�8R0�CH- YDMAXvNS_�1�1A'MOD�2AI� o �2A� (1APWD  � LA �0��ND)ATRYsFD�ELA�C2@�'`AE�RSI�1A�'RO.�ICLK�HMt0�'ί XML+ \3SG�FRM�3T� XO�U�3Z G_��COAPc1V�3Q�'C�2-5R_AU�� � �XRN1oUPDXP�COU�!SFO 3 
$V~W8o�@YACC�H�Q�SNAE$UMMY�1�W2v$DM�	�  $DISܤ�SMB�
 7T �	BCl@DC1I2AI&P6�EXPS�!�PA�R� `RANe@ � �UCL�� <(C�0�S�PTM
U� PWR8�-hCf ��Po� l5��!�"%�7Y�P�% 0�f�R�0�eP� _DL�V�De�QNIFF>� � �$?ܢBs_ST�$�: GG�$\qSv�PP̢$�@yvBUFF�&RP�q��3�IFI��>XPOSAV�dND�!\3� z��0WERUE%��EOWN��AEa0�dDe  )po�!3 
j�hX_!`�#?Z_INDE,CQ��O�pE�dUR`�D����   �t �!pMON����D���HOU�#EyA��ǁ��ǁ���LOCA� Y$�N�0H_HE���PI"/  d	`ARP�&�1�q��W_~ EwDEFS�;FA�D�01#�GHO_� �R�2P$`ށS�TEL	$# P K  !�0KWO�` Yp�PE� �LV�k�2�K IcCE����$V�  ����J��
��
���`S$Q��  �1N�$'0 	�
���F�����E��>��$� 3&������v�W��� &���!򑼯�����&������*�$;�>�ܣ�_V`&��E�l�~������� ƿؿ���� �2�פ.� _FLUp �1�W �������!�Ыnx&�2Ы*�{SHE`D 1&�Ed P���;��� ���,���P��t�7� ��[ߩ��ߑ��ߵ�� ��:���^�!�3��W� ��{���� �����6� ��Z��~�A���e��� �������� ��D P+y�a��� �
�.�d' �K�o���/ �*/�N//r/5/k/��/�/�/�/�/ԧPP�P_L�A1W�x/!1.+20�/�&�*51;?�&2551.s52?�#�C�)320?B>�0V?h?z?�?�63�?B>@�?�?�?O�64 OB>�@FOXOjO|O�65�OB>P�O�O�O�O�66_B>�P`6_H_Z_l_F�RC:�����(������{�?� Q� �/�^<"oWoio<o�o�o�o�o�o�o�(P�o) ;�o_q��T����^��)F�'���
ZDT Status�6�x�������'}iRC�onnect: �irc��//alertT������ ��f�K�]�o�������ʷ!3�P�b<��� �������(�:�L��^�p���������C�$�$c962b37�a-1ac0-e�b2a-f1c7�-8c6eb57�5d8f8  ( :��^�/�A�S�e��%)tQ��h�b�������P���`d,$&�㿚�1ѿ��� 2��?�h�Oό�sϰ� �ϩ�����
����@��'�d�K߸ ����5�PDM_�Q	�;2SMB 
 5e�3^߸_������ I�[�^��KB��_CLN�T 39+�4���n��\��� ������������C� "�g�y�X�����������.SMTP_CT�RL D��P% ��&�t��U��D�}h����NIFOF �!���"�  fr�:sniff.c�ap	frs:�diss��.dg���Ò� �Xj�������%�17�0�Q0�_��^)�����0�S��USTOM �����$` |�$�TTCPIP�Q����eb �EL325a��H!T:t/�rj3_tpd� 0P!K�CL|/put�otu��(!�CRT�/P�-?!CONS#?��!ib_smo	n+<��