��  ]i�A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ����SG_PPD�_T   � �$*ENB � $MANCM�P:F_PRES�S> $BR { ]TIMEf ]jSCLfW`
Wo	W}A_� p� ~4�* PAR�AM-   o$INI} ALs � $FFOFF�_ITP��4�& * CFG-�D $NUM_���PX6CUS�TOM�DE| H{APs $DF	�GMAX&S_EXTRA_LO��[$dNGtp�REA��SWT�CHKO_PLS�WIDTH> $�!� TMOD�D�IoOUT�US�EPROF4PM�O>!_WTLIl3�HO!MSz��TRUNCER:�F�_CH���ASSERTM��O_FCTHReS��)SE��pT:)IO�- � 
�T�AT_�^ EXI�NtPV�jEX���(� �'�!�' � �(��'�"�&]&F ~- | $�!__IOTY5sID[!4SLO@<[ 3TRCP�?0�D u!*5DINAC�KX=��GAIN�} \$S�T �\ +$C�OMMEN��$WELDSTH�ICKNVPUS�H_D 9#GUNgSAG�"<!OF	0�OUC��F�T�A:#�3== YNC��6BIER3BA�CC4CEL_R+AT;4R~ S*GPD9E�0OPN�8rBD pD,FpC9E�0_90� @ AWAY*G�B9E�To�1q x$= TR�OKE_L�B$_MOTIOt@Y:2�PEE�+AWR�3_9@_�l5U�B�6P� U�aPAT�H8V^V?�XNU�2OA_S+ G@Y�MaVD�PP@>'CRE�S02Y�S��P�8_[�VY�YZ~�8THKTBL- � � �9�:4��$$CL#   ����2a��z��'`VERS P�/h  �1N�$1 3� Ph c �v��B��� �a �i�a���o�o�o�o�o �o�o{~oLr \n���2�� ���"�H�n�X�j� �������ď֏��� ��D���H�Z����� ������ҟ�r����  ���P�b��������� 8��ԯ���(�:� L�^���������̿� ܿ� ��$ϲ�<�N� `�6ϐϢ��������� x�*��&�D�V�h�z� �ߞ���>������2� �.�@�R�d���|�� ��v������.��*� ��j�T�f��������� ����~�Lr \n���2�� ��"HnXj �������� //D/�H/Z/�/�/ �/�/�/�/�/r/�/?  ?�/P?b?�?�?�?�? 8?�?�?�?OO(O:O LO^O�O�?�O�O�O�O �O�O __$_�O<_N_ `_6_�_�_�_�_�_�_ x_*oo&oDoVohozo �o�o�o>o�o�o2 .@Rd�o|� �v���.��*� �j�T�f��������� ̏ޏ�~���L�r� \�n�������2���Ο �����"�H�n�X�j� ��������į֯��� ��D���H�Z����� ������ҿ�r����  ���P�bψϮϘϪ� 8���������(�:� L�^߄��ψߚ����� ���� ��$��<�N� `�6����������� x�*��&�D�V�h�z� ������>�����2 .@Rd��|� �v��.* �jTf���� ��/~//L/r/ \/n/�/�/�/2/�/�/ �/�/?"?H?n?X?j? �/�?�?�?�?�?�?�? OODO�?HOZO�O�O �O�O�O�O�OrO�O_  _�OP_b_�_�_�_�_ 8_�_�_�_oo(o:o Lo^o�o�_�o�o�o�o �o�o $�o<N `6������ x*��&�D�V�h�z� ����ď>�ȏڏ�2� �.�@�R�d��|��� ��v�П��.��*� ��j�T�f��������� ̯ޯ�~���L�r� \�n�������2���ο ࿶��"�H�n�X�j� ���ϔϦ��������� ��D߾�H�Zߌ߲� �߮�������r����  ���P�b����� 8���������(�:� L�^������������ ���� $��<N `6������ x*&DVhz ���>��/2/ /./@/R/d/�|/�/ �/v/�/�/?.??*? �/j?T?f?�?�?�?�? �?�?O~?OOLOrO \OnO�O�O�O2O�O�O �O�O_"_H_n_X_j_ �O�_�_�_�_�_�_�_ ooDo�_HoZo�o�o �o�o�o�o�oro�o  �oPb���� 8�����(�:� L�^��������̏� ܏� ��$���<�N� `�6�����ȟ�؟� x�*��&�D�V�h�z� ����į>�ȯگ�2� �.�@�R�d��|��� ��v�п��.��*� ��j�T�fτϖϨϺ� �����~���L�r� \�n߀ߒߤ�2߼��� �߶��"�H�n�X�j� �ߪ����������� ��D���H�Z����� ����������r���  ��Pb���� 8���(: L^������ �� //$/�</N/ `/6/�/�/�/�/�/�/ x/*??&?D?V?h?z? �?�?�?>?�?�?O2O O.O@OROdO�?|O�O �OvO�O�O_.__*_ �Oj_T_f_�_�_�_�_ �_�_o~_ooLoro \ono�o�o�o2o�o�o �o�o"HnXj �o������� ��D��H�Z����� ������ҏ�r����  ���P�b��������� 8��ԟ���(�:� L�^���������̯� ܯ� ��$���<�N� `�6�����ȿ�ؿ� x�*��&�D�V�h�z� �Ϟ���>������2� �.�@�R�d���|ߎ� ��v������.��*� ��j�T�f����� �����~���L�r� \�n�������2����� ����"HnXj�t�$SGPPD�2 3 ����� c ������� 	-?��Wi{ Q���	/�/� E///A/_/q/�/�/�/ �/�/Y/�/�/'?M?7? I?[?m???�?�?�? �?O�?#OIO3OEO�? �OoO�O�O�O�O�O_ �O_�O#_5_g_�_w_ �_�_�_�_M_�_�_�_ �_So=oco�oso�oo �o�o�o�o�oO 9_�ocu��� ������)�;� ���}���ɏ��ŏS� ����1�C�U��� y������������ 	��-�?�͟W�i�{� Q�ӯ���	����� E�/�A�_�q�����Ͽ ��߿Y����'�M�7� I�[�m��ϗϩϻ� �����#�I�3�E��� ��o߁ߟ߱������ ����#�5�g��w� �����M������� ��S�=�c���s���� ����������O 9_��cu��� �����); �}����S /�//1/C/U/�/ y/�//�/�/�/?�/ 	??-???�/W?i?{? Q?�?�?�?	O�?O�? EO/OAO_OqO�O�O�O �O�OYO�O�O'_M_7_ I_[_m___�_�_�_ �_o�_#oIo3oEo�_ �ooo�o�o�o�o�o �o�o#5g�w ����M��� �S�=�c���s���� ŏ����ߏ���O� 9�_�ُc�u���͟�� ɟ۟������)�;� ���}���ɯ��ůS� ����1�C�U��� y������������ 	��-�?�ͿW�i�{� Q��Ͻ���	���ߓ� E�/�A�_�q߃ߕ��� ����Y�����'�M�7� I�[�m������ �����#�I�3�E��� ��o����������� ����#5g�w ����M��� �S=c�s� �����//O/ 9/_/�c/u/�/�/�/ �/�/�/�/�/?)?;? ?�?}?�?�?�?�?S? O�?OO1OCOUO�O yO�OO�O�O�O_�O 	__-_?_�OW_i_{_ Q_�_�_�_	o�_o�_ Eo/oAo_oqo�o�o�o �o�oYo�o�o'M7 I[m��� ���#�I�3�E�� ��o�������ÏՏ� �����#�5�g���w� ��������M�ן��� џS�=�c���s���� ů����߯���O� 9�_�ٯc�u���Ϳ�� ɿۿ������)�;� ϓ�}ϣ��ϳ���S� �����1�C�Uߏ� yߟ�ߣߵ������ 	��-�?���W�i�{� Q������	������ E�/�A�_�q������� ����Y�����'M7 I[m��� ��#I3E� �o�����/ �/�#/5/g/�/w/ �/�/�/�/M/�/�/�/ �/S?=?c?�?s?�?? �?�?�?�?�?OOOO 9O_O�?cOuO�O�O�O �O�O�O�O�O_)_;_ _�_}_�_�_�_�_S_ o�_oo1oCoUo�o yo�oo�o�o�o�o 	-?�oWi{ Q���	���� E�/�A�_�q�����Ϗ ��ߏY����'�M�7� I�[�m��������� �����#�I�3�E�ӟ ��o�������ïկ� �����#�5�g���w� ��������M�׿��� ѿS�=�cω�sυ�� �ϯ���������O� 9�_���c�uߧ��߷� �������ߍ��)�;� ��}�������S� �����1�C�U��� y������������ 	-?��Wi{ Q���	�� E/A_q��� ��Y��'/M/7/ I/[/m///�/�/�/ �/?�/#?I?3?E?�/ �?o?�?�?�?�?�?O �?O�?#O5OgO�OwO �O�O�O�OMO�O�O�O �OS_=_c_�_s_�__ �_�_�_�_�_ooOo 9o_o�_couo�o�o�o �o�o�o�o�o); �}����S ����1�C�U��� y������������ 	��-�?�͏W�i�{� Q�ӟ���	����� E�/�A�_�q�����ϯ���߯�$SGPP�D3 3 ����$� c �Y����C�i� S�e�w�����M���ſ ׿��/��?�e�O�a� ￡ϋϝϻ������� +��;ߵ�?�Q߃ߩ� �ߥ߷�����i���� ���o�Y����� /�����������1� k�U�{���������� ������	��3E W-������ o!;M_q ���5��/)/ /%/7/I/[/�s/�/ �/m/�/�/�/%??!? �/a?K?]?{?�?�?�? �?�?�?u?�?OCOiO SOeOwO�O�O)O�O�O �O�O/__?_e_O_a_ �O�_�_�_�_�_�_�_ +oo;o�_?oQo�o�o �o�o�o�o�oio�o �ooY��� /������1� k�U�{�����Ï� ӏ���	����3�E� W�-��������ϟ� o�!���;�M�_�q� ������5���ѯ�)� �%�7�I�[��s��� ��m��ٿ��%��!� ��a�K�]�{ύϟϱ� ������u����C�i� S�e�w߉ߛ�)߳��� �߭�/��?�e�O�a� �ߡ���������� +��;���?�Q����� ����������i��� ��oY��� /����1 kU{���� ���	//�3/E/ W/-/�/�/�/�/�/�/ o/!???;?M?_?q? �?�?�?5?�?�?O)O O%O7OIO[O�?sO�O �OmO�O�O�O%__!_ �Oa_K_]_{_�_�_�_ �_�_�_u_�_oCoio Soeowo�o�o)o�o�o �o�o/?eOa �o������� +��;��?�Q����� ������ɏۏi��� ��o�Y�������� /��˟ݟ����1� k�U�{������ï� ӯ���	����3�E� W�-��������Ͽ� o�!���;�M�_�q� �ϕϻ�5Ͽ����)� �%�7�I�[���s߅� ��m�������%��!� ��a�K�]�{���� ������u����C�i� S�e�w�����)����� ����/?eOa ��������� +;�?Q�� �����i�/ /�o/Y//�/�/�/ //�/�/�/�/??1? k?U?{?�/?�?�?�? �?�?�?	OO�?3OEO WO-O�O�O�O�O�O�O oO!___;_M___q_ �_�_�_5_�_�_o)o o%o7oIo[o�_so�o �omo�o�o�o%! �oaK]{��� ���u��C�i� S�e�w�����)���ŏ ׏��/��?�e�O�a� �������͟ߟ� +��;���?�Q����� ������ɯۯi��� ��o�Y�������� /��˿ݿ����1� k�U�{���ϑ����� ������	�ߩ�3�E� W�-߯ߙ߿������� o�!���;�M�_�q� ����5�����)� �%�7�I�[���s��� ��m�������%! ��aK]{��� ���u�Ci Sew��)�� ��///?/e/O/a/ ��/�/�/�/�/�/�/ +??;?�/??Q?�?�? �?�?�?�?�?i?�?O O�?oOYOO�O�O�O /O�O�O�O�O__1_ k_U_{_�O_�_�_�_ �_�_�_	oo�_3oEo Wo-o�o�o�o�o�o�o oo!;M_q ���5���)� �%�7�I�[��s��� ��m��ُ��%��!� ��a�K�]�{������� �՟��u����C�i� S�e�w�����)���ů ׯ��/��?�e�O�a� ﯡ�������Ϳ߿� +��;ϵ�?�Qσϩ� �ϥϷ�����i���� ���o�Y�ߥߏߡ� /�����������1� k�U�{��������� ������	����3�E� W�-������������� o�!;M_q ���5��) %7I[�s� �m���%//!/ �a/K/]/{/�/�/�/ �/�/�/u/�/?C?i? S?e?w?�?�?)?�?�? �?�?/OO?OeOOOaO �?�O�O�O�O�O�O�O�+__;_�$SGP�PDCFG �����Q�  u P��P  �_P�O_]R�_ZU�Q�S�@\S�WX2�BH��VuTIO1 3��[c �]UQ_ YY)oGo9oKo}ooo �o�o�o�o�o�o�o�o %UCYk�� �������3� Q�C�i�c�u������� Տ���%��A�_� Q�w�������ǟ��� ���7�)�O�i�[� ��������ٯ˯t�� ��'�E�7�]�{�m��� ����ɿ�ٿ��� 1�O�A�Wω�{ύϟ� �Ͽ��������1�/� A�g�a�sߝߛ߭��� ����	���?�]�O� u����������� ���5�'�M�g�Y��� ������������	�� %C5[yk� �����R M?i�y��� ����)//-/?/ e/_/�/�/�/�/�/�/ �/???=?;?M?s? �?�?�?�?�?�?�?�? O3O%OKOeOWO�O�O �O�O�O�O�O_�O#_ A_3_Y_w_i_�_�_�_ �_�_�_�_oo�_Ko =ogo�owo�o�o�o�o �o�o	'+]O q������� ��5�#�9�K�q�o� ��������ݏۏ�� 1�#�I�C�U������ ��ӟş����!�?� 1�W�u�g�������ï �ӯ���	�/�I�;� e���u�������T�� ݿ�%��=�[�Mϒ� ��ϩ��Ϲ������� �/�!�7�i�[�m�� �ߟ����������� !�G�A�S�}�{��� �����������=�/� U�s�e����������� ����-G9c �s������ #;YK�� }������2/ -//I/g/Y/k/�/�/ �/�/�/�/	?�/?? E???u?c?y?�?�?�? �?�?�?�?OO-OSO qOcO�O�O�O�O�O�O �O__+_E_7_a__ q_�_�_�_�_�_�_o !oo9oWoIooo�o{o �o�o�o�o�o�o�o+ GeW}��� ������=�/� Q�o�a�w��������� �ߏ���+�Q�O� a�����������͟� ��)�#�5�_�}�o� ������˯�ׯ�� �7�U�G�m���y��� ����ٿ����)�� E�c�U�{ϙϋ�4��� ��������;�-�r� m�_߉ߧߙ߫����� �����I�;�M�_� ������������ �'�!�3�]�[�m��� ������������ 5SEk�w�� ����'C aSy����� �/�/9/+/�k/ ]/�/�/�/�/�/�/? ?�/)?G?9?K?}?o? �?�?�?�?�?�?�?�? %OOUOCOYOkO�O�O �O�O�O�O�O�O_3_ Q_C_i_c_u_�_�_�_ �_�_�_o%ooAo_o Qowo�o�o�o�o�o�o �o7)Oi[ ������t� �'�E�7�]�{�m��� ����ɏ�ُ��� 1�O�A�W���{����� ş��������1�/� A�g�a�s�������ӯ ��	���?�]�O� u�������ſ����� ��5�'�M�g�Yσ� �ϓϹ�������	��� %�C�5�[�y�k�߫� ������������R� M�?�i��y���� ��������)��-�?� e�_������������� ��=;Ms �������� 3%KeW�� �����/�#/ A/3/Y/w/i/�/�/�/ �/�/�/�/??�/K? =?g?�?w?�?�?�?�;��$SGPPDI�O2 3����A c ��?�?#OAO3O YOwOiOT?�O�O�O�O �O�O__P_K_=_g_ �_w_�_�_�_�_�_�_ �_'oo+o=oco]o�o �o�o�o�o�o�o�o ;9Kq��� ������1�#� I�c�U��������ӏ ŏ����!�?�1�W� u�g�������ß�ӟ ���	���I�;�e��� u���������ݯ� %��)�[�M�o���� ��ǿ��˿ݿ���3� !�7�I�o�m�ϥϟ� ���������/�!�G� A�S�}ߛߍ߳����� ������=�/�U�s� e������������ ��-�G�9�c���s� ������R�����# ;YK��}� �����- 5gYk}��� ���///E/?/ Q/{/y/�/�/�/�/�/ �/�/?;?-?S?q?c? �?�?�?�?�?�?�?O O+OEO7OaOOqO�O �O�O�O�O�O_!__ 9_W_I_�O�_{_�_�_ �_�_�_�_0o+ooGo eoWoio�o�o�o�o�o �o�oC=s aw������ ���+�Q�o�a��� ������ۏ͏��� )�C�5�_�}�o����� ��˟�ן���7� U�G�m���y������� ٯ��鯒�)��E�c� U�{�����п˿��� ���	�;�-�O�m�_� uϧϙϫϽ������ ��)�O�M�_߅�� �߻߹�������'� !�3�]�{�m���� ����������5�S� E�k���w��������� ����'CaS y��2��� �9+pk]� ������/� /G/9/K/]/�/}/�/ �/�/�/�/�/�/%?? 1?[?Y?k?�?�?�?�? �?�?�?OO3OQOCO iO�OuO�O�O�O�O�O �O_%__A___Q_w_ �_�_�_�_�_�_o�_ o7o)o�_io[o�o�o �o�o�o�o�o' E7I{m��� �����#��S� A�W�i�������ŏ�� я�����1�O�A�g� a�s�������ӟ�� 	�#��?�]�O�u��� ����ů������� 5�'�M�g�Y������� ��׿ɿr�	���%�C� 5�[�y�kϰϫϝ��� ��������/�M�?� U߇�yߋߝ��߽��� ����	�/�-�?�e�_� q����������� ��=�[�M�s����� ������������3 %KeW���� ����#A3 Ywi���� ��//P/K/=/g/ �/w/�/�/�/�/�/�/ �/'??+?=?c?]?�? �?�?�?�?�?�?O�? O;O9OKOqO�O�O�O �O�O�O�O�O_1_#_ I_c_U__�_�_�_�_ �_�_o�_!o?o1oWo uogo�o�o�o�o�o�o �o	�oI;e� u������� %��)�[�M�o���� ��Ǐ��ˏݏ���3� !�7�I�o�m������ ��ٟ۟��/�!�G� A�S�}�������ѯï �����=�/�U�s� e���������߿ѿ�� ��-�G�9�cρ�s� �Ϸϩ�R������#� �;�Y�Kߐߋ�}ߧ� �߷��������-�� 5�g�Y�k�}����� ���������E�?� Q�{�y����������� ����;-Sqc ������� +E7aq������$SGP�PDIO3 3����!? c ��� !/?/1/W/u/g/R�/ �/�/�/�/�/?	?N? I?;?e?�?u?�?�?�? �?�?�?�?%OO)O;O aO[O�OO�O�O�O�O �O_�O_9_7_I_o_ �__�_�_�_�_�_�_ o/o!oGoaoSo}o�o �o�o�o�o�o�o =/Use��� �������G� 9�c���s�������� �ۏ�#��'�Y�K� m���}���ş��ɟ۟ ���1��5�G�m�k� }�������ٯׯ�� -��E�?�Q�{����� ��Ͽ������;� -�S�q�cωϣϕϿ� ��������+�E�7� a��qߗߵߧ�P��� ���!��9�W�I�� ��{����������� �+��3�e�W�i�{� ������������ C=Oyw�� �����9+ Qoa����� ��//)/C/5/_/ }/o/�/�/�/�/�/�/ ???7?U?G?�/�? y?�?�?�?�?�?�?.O )OOEOcOUOgO�O�O �O�O�O�O_�O	__ A_;_q___u_�_�_�_ �_�_�_�_oo)oOo mo_o�oo�o�o�o�o �o'A3]{ m������� ��5�S�E�k���w� ������׏��珐�'� �C�a�S�y�����Ο ɟ�������9�+� M�k�]�s��������� �ۯ����'�M�K� ]���}�������ɿ� ���%��1�[�y�k� �ϯϡ���������� �3�Q�C�i߃�uߟ� �߯��������%�� A�_�Q�w���0��� ��������7�)�n� i�[������������� ����E7I[ �{������ �#/YWi� ������// 1/O/A/g/�/s/�/�/ �/�/�/�/	?#???? ]?O?u?�?�?�?�?�? �?�?�?O5O'O�?gO YO�O�O�O�O�O�O_ 	_�O%_C_5_G_y_k_ �_�_�_�_�_�_�_�_ !ooQo?oUogo�o�o �o�o�o�o�o�o	/ M?e_q��� ����!��=�[� M�s�������Ï��ߏ ����3�%�K�e�W� ��������՟ǟp�� ��#�A�3�Y�w�i��� ����ů�կ��� -�K�=�S���w����� �����߿���-�+� =�c�]�oϙϗϩ��� ��������;�Y�K� qߏ߁ߧ��߳����� ���1�#�I�c�U�� ������������� !�?�1�W�u�g���� ����������	N I;e�u��� ����%); a[����� �/�/9/7/I/o/ �//�/�/�/�/�/�/ ?/?!?G?a?S?}?�? �?�?�?�?�?O�?O =O/OUOsOeO�O�O�O �O�O�O�O__�OG_ 9_c_�_s_�_�_�_�_ �_�_o#oo'oYoKo mo�o}o�o�o�o�o�o �o15Gmk }������� -��E�?�Q�{����� ��Ϗ������;� -�S�q�c��������� ݟϟ����+�E�7� a��q�������P�� ٯ�!��9�W�I��� ��{���ÿ��ǿ��� �+��3�e�W�i�{� �ϛ��Ͽ������� �C�=�O�y�w߉߯� �߿��������9�+� Q�o�a������� ������)�C�5�_��}�o����������$�SGPPDSET�1 ���^����wB?���BH���2 �� 23�CUgSCH1 �1c �
�Producti{on��C�����@@��A�  ���� d dB � ��	� 4�� �6��� ��j����&8J\�
���~��������
��/0/B/�T/f/x/�/�/�
�o߾/�/�/�/??*?<?�
���^?p?�?��?�?�?�?�?�
���?O"O4OFOXOjO|O�
�tݞO�O�O��O�O�O
__�
���>_P_b_t_�_�_�_�_�
�"��_�_o�o&o8oJo\o�
�y�~o�o�o�o�o�o�o<�o�	Dhb0�BTfx���z������8*�<��z�\^�p����������ʏ܏�z |� �2�D�V�h�z��|f����ԟ`���
���z� O�a�s����������{$m`ޯ���&�p8�J�\��z*�~� ������ƿؿ����z/�Z�0�B�T�f�xϊϜϮz5\?���������(�:߬|;T^�p߂ߔߦ߸����߮z@�����"��4�F�X�j�|�zFr^�����������
���zL�ON�`�r���p�������|Q�X�� ��&8J\n
W<_��������|] R0B�Tfx��n
b�׾���//*/</n
hwL^/p/�/@�/�/�/�/�/n
n|o ? ?2?D?V?h?z?�|s�V�?�?�?�?�?p�?
OOn
yy�>O PObOtO�O�O�O�On
%P�O�O__&_8_J_\_n
���_�_ �_�_�_�_�^�[$f"o 4oFoXojo|o�o�o�o �o�o�o�o0B Tfx����� ����,�>�P�b� t���������Ώ��� ��(�:�L�^�p��� ������ʟܟ� �� $�6�H�Z��~����� ��Ưد����� �2� D�V�h�z�����O�¿ Կ���
��.�@�R� d�vψϚϬϾ����� ����*�<�N�`�r� �ߖߨߺ�������� �&�8�J�\�n�������aForce�Check��C�������&�8�qJ�\�n�#K~� ��������������n��|�.@Rdv��l��o߾����*<n����^p������n��y��/"/�4/F/X/j/|/n�D�/�/�/�/�/�/8
??.:j�>?P?�b?t?�?�?�?�?.:��/�?OO%O7OIO[O-;*�~O�O�O@�O�O�O�O�O.:5\ ._@_R_d_v_�_�_,<@�پ_�_�_�_opo*o<o.:L�^o po�o�o�o�o�o�o.:Wt��o"4FpXj|.:b�מ �����
��.:n"�>�P�b�t���p������.:yy�ޏ ����&�8�J�\�.:�hb~�������Ɵ ؟ꟼﭯ �2�D�V� h�:�����O�¯ԯ� ��
��.�@�R�d�v� ��������п���� �*�<�N�`�rτϖ� �Ϻ���������&� 8�J�\�n߀ߒߤ߶� ���������"�4�F� X�j�|�������� ������0�B�T�f� x�����M�������� ,>�bt� ������ (:L^p��� ���� //$/6/ H/Z/l/~/�/�/�/�/ �/�/�/? ?2?D?V? h?z?�?�?�?�?�?�? �?
OO.O@OROdOvO �O�OK_�O�O�O�O_ _*_<_�_`_r_�_�_ �_�_�_�_�ooo&o 8oJo\ono�o�o�o�o��o�o�o�o�	I�nsertCapHrC��uFX�j|����uTip Dress�s#K>���&��8�J���TD New �tz��������ԏ���
Sit�PrsNwC��o�0|-�?�Q�c�u������
Resis�t Chk�r���П�����*��\�Deburr e���b�t����������ί �Auto�lib6��,�>�P��b�t�f�L�erve������¿Կ��� 
��.�@�R�d�vψ��Ϭ�~� 0�����?@��dA���0~����#�5�G�Y���AW"�� �� �߀�ߴ�������������$SGSCH2 �1������ c ��
ProductionV�����L��^��߂�����j��������"�4�F�X�����z�������������������,>Pbt� ���������8#5�����Zl�~����������//0/B/T/8f/x/���tݚ/�/��/�/�/�/??�����:?L?^?p?�?�?8�?�?���"��?�?��?O"O4OFOXO���y�zO�O�O�O�O�O8�O�O��Dh��_ 0_B_T_f_x_�_�_�V�_�_�_�_opo&o8o�Z�\Zo lo~o�o�o�o�o�o�Zx�
.@Rdv�\f����������Z� _K�]�o����������[$m`ڏ�����"�4�F�X��Z*� z�������ԟ����Z/�Z�,�>�P� b�t������Z5Xʯ�ܯ� ��$�6��\;TZ�l�~�������8ƿؿ�Z@����π�0�B�T�f�xϪZFr^�ϬϾ��������ߪZL�/J�\�n���ߒߤ߶ߨ\Q�X �������"�4�F�X�j�W8?��������8����\] R�,��>�P�b�t�����j�b�׺�������8&8j�hwLZl�~�����j�n xO
.@Rdv�\s�V�������//j�yy� :/L/^/p/�/�/�/�/j�%P�/�/�/? "?4?F?X?jꂸ_�? �?�?�?�?�?�>�; F O0OBOTOfOxO�O�O �O�O�O�O�O__,_ >_P_b_t_�_�_�_�_ �_�_�_oo(o:oLo ^opo�o�o�o�o�o�o �o $6HZl ~������� � �2�D�V��z��� ����ԏ������ .�@�R�d�v�����K� ��П�����*�<� N�`�r���������̯ ޯ���&�8�J�\� n���������ȿڿ� ���"�4�F�X�j�|���Ϡϲ�AForc�eCheck��C��������"��4�F�X�j�#K zߌߞ߰���������jڈY+�=�O�a�ps���i۵oߺ� ��������&�8�j����Z�l�~�����p������j��y��� 0BTfxj�D�������*j� :L^p����*����/!/p3/E/W/)*�z/ �/�/�/�/�/�/�/*5X�*?<?N?`?r?�?�?(@�ٺ?�?�?��?OO&O8O*L�ZOlO~O�O�O�O�O�O*Wt��O__�0_B_T_f_x_*b� ��_�_�_�_�_oo)n"�:oLo^opo��o�o�o�o*yy� �o�o�o"4FX*�hbz��� ����ϩ��.�@� R�d�6߈���K���Џ ����*�<�N�`� r���������̟ޟ� ��&�8�J�\�n��� ������ȯگ���� "�4�F�X�j�|����� ��Ŀֿ�����0� B�T�f�xϊϜϮ��� �����ϧ��,�>�P� b�t߆ߘ�I������ ����(�:���^�p� ����������� � �$�6�H�Z�l�~��� ������������  2DVhz��� ����
.@ Rdv����� ��//*/</N/`/ r/�/�/G?�/�/�/�/ ??&?8?�?\?n?�? �?�?�?�?�?�O�?O "O4OFOXOjO|O�O�O��O�O�O�O�O_�v	�InsertCa=pDRC�:_L_�^_p_�_�_�_�]Tip Dress�S#K�_�_�_o"o�4oFo�}TD New �Tvo�o�o�o�o��o�o�o
Sit�PrsNwCs�o�,>Pbt���mResist� Chk�R�� ������&�XlDeburra� �h�z�������ԏ�
Autoplib2_��(�:�L��^�p�"RH�erve��������П��� ��*�<�N�`�r��� ������̯ޯ��� &�8�J�\�n�������඿ȿڿ�!��$S�GSCH3 1������? c �&_� *�<�N�`�rτ�_c� ��������0�B�T� �xߊߜ߮������� �ߧ��,�>�P�b�t� ������������ �(�:�L�^�p����� ���������� $ 6HZl~��� ���� 2D Vhz����� ��
//./@/R/? v/�/�/�/�/�/�/�/ �??*?<?N?`?r?�? �?GO�?�?�?�?OO &O8OJO\OnO�O�O�O �O�O�O�O�O_"_4_ F_X_j_|_�_�_�_�_ �_�_�_oo0oBoTo foxo�o�o�o�o�o�o �o,>Pbt ��������� �(�:�L�^�p����� E���ʏ܏� ��$� 6��Z�l�~������� Ɵ؟���� �2�D� V�h�z�������¯ԯ ���
��.�@�R�d� v���������п��� ��*�<�N�`�rτ� �ϨϺ��������� &�8�J�\�n߀ߒ�C� �����������"�4� ��X�j�|������ �������0�B�T� f�x������������� ��,>Pbt ������� (:L^p�� ����� //$/ 6/H/Z/l/~/�/�/�/ �/�/�/�/? ?2?�? V?h?z?�?�?�?�?�? �O�?
OO.O@OROdO vO'_�O�O�O�O�O�O __*_<_N_`_r_�_ �_�_�_�_�_�_oo &o8oJo\ono�o�o�o �o�o�o�o�o"4 FXj|���� �����0�B�T� f�x���������ҏ�� ����,�>�P�b�t� %�������Ο���� �ǯ:�L�^�p����� ����ʯܯ� ��$� 6�H�Z�l�~������� ƿؿ���� �2�D� V�h�zόϞϰ����� ����
��.�@�R�d� v߈ߚ߬߾������� ��*�<�N�`�r�#� ������������ ��8�J�\�n������� ��g������"4 FXj|���� ���0BT fx������ �//,/>/P/b/t/ �/�/�/�/�/�/�/? ?(?:?L?^?p?�?�? �?�?�?�?�? OO�O 6OHOZOlO~O�O�O�O e_�O�O�O_ _2_D_ V_oz_�_�_�_�_�_ �_�_
oo.o@oRodo vo�o�o�o�o�o�o�o *<N`r� �������� &�8�J�\�n������� ��ȏڏ����"�4� F�X�j�|�������c� ֟�����0�B�T� �x���������ү� �����,�>�P�b�t� ��������ο��� �(�:�L�^�pςϔ� �ϸ������� ��$� 6�H�Z�l�~ߐߢߴ� ��������� �2�D� V�h�z�������� ����
��.�@�R� v��������������� �*<N`r� �G���� &8J\n��� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO �O�O�O�O�O�O�O�_ _(_:_L_^_p_�_�_ Eo�_�_�_�_ oo$o 6o�oZolo~o�o�o�o �o�o�o�o 2D Vhz����� ��
��.�@�R�d� v���������Џ�� ��*�<�N�`�r����������̟ޟ��$�SGTHKTBL�1 2������ 
� CalGoauge�AP ��	PartThick��ӯ������� �2�D�V�h���2 ����ѯ�m�ڿ��� �"�4�FϞ�3���� �~��ϡϳ������� ����1�