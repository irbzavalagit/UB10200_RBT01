��   X�A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ����CIPS_C�FG_T   �0 $INTE�RFACE  �$DUMMY1�B2B3B&SE�T/ @ $�MODA8 _S�IZ}OUT�DATE_FIX~�CSI_VRC �  4��$$CLASS ? �������O��O� VERS�ION�  1N�$'1 �O� �m �r �
���  . 0-@