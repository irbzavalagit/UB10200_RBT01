��   (�A��*SYST�EM*��V9.3�0126 2/�12/2021 A 	  ����PASSNA�ME_T   �0 $+ �$'WORD � ? LEVEL � $TI- OUTT4&F/�� $SE�TUPJPROG�RAMJINST�ALLJY  $CURR_OަUSER�NU�M�STSTOP�_TPCHG �V LOG_P NT��N�  6 C�OUNT_DOW�N�$ENB_�PCMPWD� �$DV_� IN�� $C� CR5E��A RM9� =T9DIAG9(|�LVCHK >FULLM/��YXT�CNTD��MENU�A�UTO+�FG_wDSP�RLS��U�BURYBA�N��GI�eE�NC/  ~CRYPTE�  �4��$$CL(   ���[!�� d �P V� IONX(�  1N��$DCS_CO�D?���_%� � Ɋ'_� �.W��(S  Z*�� $\ �&�A91�"[!�	 
 �$��011��  0b!;��6?k?Z?�? ~?�?�?�?�?�?�?O�OCO2OgO�#SUP
�  :�?$?�#F��KWM�O�� � \Q��_ �0�� V�[_t&��j��.4hOp_��.W,_�� �V�U�YqILUGH� 1[) � �)�_oo/o AoSoeowo�o�o�o�o �o�'�_�o#5G Yk}����� �o���1�C�U�g� y���������ӏ�� 	��-�?�Q�c�u��� ������ϟ����� )�;�M�_�q������� ��˯ݯ���%�7� I�[�m��������ǿ ٿ����!�3�E�W� i�{ύϟϱ������� ����/�A�S�e�w� �ߛ߭߿�������� �+�=�O�a�s��� ��������� ��'� 9�K�]�o��������� ���������#5G Yk}����� ���%