��   G-�A��*SYST�EM*��V9.3�0126 2/�12/2021 A   ����SG_DST�_T   � �$COMMEN�T $*G�UN  BR�B= L R, ERM�TYPJ ZAC�CeAP]
u MO>|SPEEDpm�EQ_ENBJ `�G� S� SP���PUSH* JL�IN)J4�$�$CLASS  �������C���C� VERSI�ON� � 1N�$SG�* 1 1 C� c <
2m�mGunOpen6��?�U d_^6��@@mA u��
4Jp�_q�
6�����
8�X!��'
10J��E#/%/7 5;)wK/]/�2v+H/�/|3v+��/�/}v*B�/?�*;p9?K?�*;�/�?0(v!/6ȱ?�?1&�"�/6�/�?0')2?%C )O;O1&e2[F8?vO0'��2[F4�O�O�&�:CaH�O�O�&JC\_�+_�&VKt?f_�'�K��_�_�&�K��_�_�&
[�	oo�&F[�?Vo l/B&{�o�oPw-�o �o/e�-�o�k(@7I5:*71s��7�{�P��9 �{4�0'9"�9'�9� 3$%rIc�u��eS�cA ����3$�r�Iۏ�3$ ��I�)��$R�QS� e��$��SQ�����%ˊ �ڟ�'��P���$ B�`C�U��$~�D`� ���$��$�ʯ�/�g�o 
� v4�F�\2sp� ���ns������� ����$�6�4$S��� n�HS��Ϯ�PD���� �όDˎ�&��D�P� b�TC��ߞ�@T��� ��|T����T��@� R��T3�|��0do��� ��ld������#.�� >��jw(@o���K�x 71������P���� �ΐPs1#5��`� _q;ݯ1�1��w�B�	�����1�1%��B܁Oa@+�'A'A��g�� ����d@cA//��q#?/Q/���A{/D�/W�*�#�/�/��6�o�/��	Tip? Dress"3�裱0?B?
U0Chn/gFix��`e?w?��<Mov�?�?��U�serCustom[��?�?O%?'O9O KO]OoO�O�O�O�O�O �O�O�O_#_5_G_Y_ k_}_�_�_�_�_�_�_ �_oo1oCoUogoyo �o�o�o�o�o�o�o	�-?~Re
@verr]o�����{g��v���F�(����$SGDS�T2 1 �������c i<k�#�eb�?��� �i�������₯��� �֋�����K�֋�� [�'�9���#�/�c�u� ��"�k��������ן ��$ƛ��%���"� ��O�a���z�X ���� ��z��֯Ƒ��� �C/�L�N�|/�;! {��������ƿ��� ����3��  /�A� o��<�k�}ϫ��į �����������#%�� � �1�_%��,�[�m� �%�� ��߼������ 3ǝ�!�_%�K�]� τ�������5��������7��X �����9����J���3�w� ��u�o�������+- ��)��+=�� e�#�gy����g�� ������������* 8�*��V�Wi�� �XГ�7����� �7�
t�/����� Z/p�.��/�/����/ �/����/?���8? J?H�*�t?�?�����/ �?`����?�?����(O :OܴdOvO�W�O �OTē�O�O���_ *_��T_f_�G�_ �_Dԃ�_�_�Կo o���DoVo8�~[�? �oX?��x��o�o�>d  ���o�>h�kq7I NT7�s�ONX��q ���M�1�1���MB�Y�'�9�]���c�u�?]B�у����@{]w�w�ۏ폷^I� �)��^��'S�e�/n������knd �˟Dݟ�n*9���!��h�G�M�#�	Tip? Dressr���!����
��Chn/gFix�"`��ǯ�٬Mov����U�serCustoms�9�K�]�o����� ����ɿۿ����#� 5�G�Y�k�}Ϗϡϳ� ����������1�C� U�g�yߋߝ߯����� ����	��-�?�Q�c�u��!�Re��ve�������������+�=�O�a�s�!���$SGDST3 �1 �����;K�c <g��� ��a���);M _q������ �%7I[m ������� /!/3/E/W/i/{/�/ �/�/�/�/�/�/?? /?A?S?e?w?�?�?�? �?�?�?�?OO+O=O OOaOsO�O�O�O�O�O �O�O__'_9_K_]_ o_�_�_�_�_�_�_�_ �_o#o5oGoYoko}o �o�o�o�o�o�o�o 1CUgy�� �����	��-� ?�Q�c�u��������� Ϗ����)�;�M� _�q���������˟ݟ ���%�7�I�[�m� �������ǯٯ��� �!�3�E�W�i�{��� ����ÿտ����� /�A�S�e�wωϛϭ� ����������+�=� O�a�s߅ߗߩ߻��� ������'�9�K�]� o����������� ���#�5�G�Y�k�}� �������������� 1CUgy�� �����	- ?Qcu���� ���//)/;/M/ _/q/�/�/�/�/�/�/ �/??%?7?I?[?m? ?�?�?�?�?�?�?�? O!O3OEOWOiO{O�O �O�O�O�O�O�O__ /_A_S_e_w_�_�_�_ �_�_�_�_oo+o=o Ooaoso�o�o�o�o�o