��   ��A��*SYST�EM*��V9.3�0126 2/�12/2021 A 	  ����DRYRUN�_T  4 �$'ENB � $NUM_P�ORTA ESU�@$STATE� P TCOL_���PMPMCmGRP_MASKZ}E� OTIONN�LOG_INFO�NiAVcFLTR_EMPTYd $PROD__ �L �ESTOP_�DSBLAPOW�_RECOVAO{PR�SAW_� �G %$IN�IT	RESUM�E_TYPEND�IST_DIFF>A $ORN41p� d =R�4&�J_  4 �$(F3IDXX��_ICIg�MIX_BG-<y
_NAMc gMODc_USd~�IFY_TI�� �MKR-�  $LIN�c   "_S�IZc�� �. �h $USE_FLC 3!�:&iF*SIMA7#Q�C#QBn'SCAN��AX�+IN�*I���_COUNrR�O( ��!_TMR�_VA�g# h>�ia �'` ����1�+WAR��$�H�!�#Nf3CH�PE�$,O�!PR�'Ioq7�iOqfOoAT�H- P $ENABL+��0BTf�$$�CLASS  O���A��5��=5�0VERS�G�  1�N�6/ E+5�������-@B]F@AbE��%A �O���O�O����3EvI2>K �O _/_A_S_e_w_�_�_ �_�_�_�_�_oo+o��O)W?"HI@ ��lj@|o�or�i�� � 2>I�  4%B�GMAI@�o���_AR�;��aAP�P1�o�o_AoAt2�%&8|3YZ8|4���8|B��<x6 ��8v)�V���c$"P+ �ktK-@����bA��X_AA-@vN ڏ����"�4�F�X� j�|���������bFoA ǁoA���
��.�@� R�d�v���������Я�DZM�_E�cC!2�lǏ1�C�U�g� y���������ӿ��� 	�Ɯ#�<�N�`�rτ� �ϨϺ��������� �8�J�\�n߀ߒߤ� �����������"�-� F�X�j�|������ ��������)�;�T� f�x������������� ��,7�Pbt ������� (:E^p�� ����� //$/ 6/ASl/~/�/�/�/ �/�/�/�/? ?2?D? Ch�4�0��{?@